magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect 0 0 856 1214
<< pmoslvt >>
rect 204 102 274 1112
rect 330 102 400 1112
rect 456 102 526 1112
rect 582 102 652 1112
<< pdiff >>
rect 148 1100 204 1112
rect 148 1066 159 1100
rect 193 1066 204 1100
rect 148 1032 204 1066
rect 148 998 159 1032
rect 193 998 204 1032
rect 148 964 204 998
rect 148 930 159 964
rect 193 930 204 964
rect 148 896 204 930
rect 148 862 159 896
rect 193 862 204 896
rect 148 828 204 862
rect 148 794 159 828
rect 193 794 204 828
rect 148 760 204 794
rect 148 726 159 760
rect 193 726 204 760
rect 148 692 204 726
rect 148 658 159 692
rect 193 658 204 692
rect 148 624 204 658
rect 148 590 159 624
rect 193 590 204 624
rect 148 556 204 590
rect 148 522 159 556
rect 193 522 204 556
rect 148 488 204 522
rect 148 454 159 488
rect 193 454 204 488
rect 148 420 204 454
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 274 1100 330 1112
rect 274 1066 285 1100
rect 319 1066 330 1100
rect 274 1032 330 1066
rect 274 998 285 1032
rect 319 998 330 1032
rect 274 964 330 998
rect 274 930 285 964
rect 319 930 330 964
rect 274 896 330 930
rect 274 862 285 896
rect 319 862 330 896
rect 274 828 330 862
rect 274 794 285 828
rect 319 794 330 828
rect 274 760 330 794
rect 274 726 285 760
rect 319 726 330 760
rect 274 692 330 726
rect 274 658 285 692
rect 319 658 330 692
rect 274 624 330 658
rect 274 590 285 624
rect 319 590 330 624
rect 274 556 330 590
rect 274 522 285 556
rect 319 522 330 556
rect 274 488 330 522
rect 274 454 285 488
rect 319 454 330 488
rect 274 420 330 454
rect 274 386 285 420
rect 319 386 330 420
rect 274 352 330 386
rect 274 318 285 352
rect 319 318 330 352
rect 274 284 330 318
rect 274 250 285 284
rect 319 250 330 284
rect 274 216 330 250
rect 274 182 285 216
rect 319 182 330 216
rect 274 148 330 182
rect 274 114 285 148
rect 319 114 330 148
rect 274 102 330 114
rect 400 1100 456 1112
rect 400 1066 411 1100
rect 445 1066 456 1100
rect 400 1032 456 1066
rect 400 998 411 1032
rect 445 998 456 1032
rect 400 964 456 998
rect 400 930 411 964
rect 445 930 456 964
rect 400 896 456 930
rect 400 862 411 896
rect 445 862 456 896
rect 400 828 456 862
rect 400 794 411 828
rect 445 794 456 828
rect 400 760 456 794
rect 400 726 411 760
rect 445 726 456 760
rect 400 692 456 726
rect 400 658 411 692
rect 445 658 456 692
rect 400 624 456 658
rect 400 590 411 624
rect 445 590 456 624
rect 400 556 456 590
rect 400 522 411 556
rect 445 522 456 556
rect 400 488 456 522
rect 400 454 411 488
rect 445 454 456 488
rect 400 420 456 454
rect 400 386 411 420
rect 445 386 456 420
rect 400 352 456 386
rect 400 318 411 352
rect 445 318 456 352
rect 400 284 456 318
rect 400 250 411 284
rect 445 250 456 284
rect 400 216 456 250
rect 400 182 411 216
rect 445 182 456 216
rect 400 148 456 182
rect 400 114 411 148
rect 445 114 456 148
rect 400 102 456 114
rect 526 1100 582 1112
rect 526 1066 537 1100
rect 571 1066 582 1100
rect 526 1032 582 1066
rect 526 998 537 1032
rect 571 998 582 1032
rect 526 964 582 998
rect 526 930 537 964
rect 571 930 582 964
rect 526 896 582 930
rect 526 862 537 896
rect 571 862 582 896
rect 526 828 582 862
rect 526 794 537 828
rect 571 794 582 828
rect 526 760 582 794
rect 526 726 537 760
rect 571 726 582 760
rect 526 692 582 726
rect 526 658 537 692
rect 571 658 582 692
rect 526 624 582 658
rect 526 590 537 624
rect 571 590 582 624
rect 526 556 582 590
rect 526 522 537 556
rect 571 522 582 556
rect 526 488 582 522
rect 526 454 537 488
rect 571 454 582 488
rect 526 420 582 454
rect 526 386 537 420
rect 571 386 582 420
rect 526 352 582 386
rect 526 318 537 352
rect 571 318 582 352
rect 526 284 582 318
rect 526 250 537 284
rect 571 250 582 284
rect 526 216 582 250
rect 526 182 537 216
rect 571 182 582 216
rect 526 148 582 182
rect 526 114 537 148
rect 571 114 582 148
rect 526 102 582 114
rect 652 1100 708 1112
rect 652 1066 663 1100
rect 697 1066 708 1100
rect 652 1032 708 1066
rect 652 998 663 1032
rect 697 998 708 1032
rect 652 964 708 998
rect 652 930 663 964
rect 697 930 708 964
rect 652 896 708 930
rect 652 862 663 896
rect 697 862 708 896
rect 652 828 708 862
rect 652 794 663 828
rect 697 794 708 828
rect 652 760 708 794
rect 652 726 663 760
rect 697 726 708 760
rect 652 692 708 726
rect 652 658 663 692
rect 697 658 708 692
rect 652 624 708 658
rect 652 590 663 624
rect 697 590 708 624
rect 652 556 708 590
rect 652 522 663 556
rect 697 522 708 556
rect 652 488 708 522
rect 652 454 663 488
rect 697 454 708 488
rect 652 420 708 454
rect 652 386 663 420
rect 697 386 708 420
rect 652 352 708 386
rect 652 318 663 352
rect 697 318 708 352
rect 652 284 708 318
rect 652 250 663 284
rect 697 250 708 284
rect 652 216 708 250
rect 652 182 663 216
rect 697 182 708 216
rect 652 148 708 182
rect 652 114 663 148
rect 697 114 708 148
rect 652 102 708 114
<< pdiffc >>
rect 159 1066 193 1100
rect 159 998 193 1032
rect 159 930 193 964
rect 159 862 193 896
rect 159 794 193 828
rect 159 726 193 760
rect 159 658 193 692
rect 159 590 193 624
rect 159 522 193 556
rect 159 454 193 488
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 285 1066 319 1100
rect 285 998 319 1032
rect 285 930 319 964
rect 285 862 319 896
rect 285 794 319 828
rect 285 726 319 760
rect 285 658 319 692
rect 285 590 319 624
rect 285 522 319 556
rect 285 454 319 488
rect 285 386 319 420
rect 285 318 319 352
rect 285 250 319 284
rect 285 182 319 216
rect 285 114 319 148
rect 411 1066 445 1100
rect 411 998 445 1032
rect 411 930 445 964
rect 411 862 445 896
rect 411 794 445 828
rect 411 726 445 760
rect 411 658 445 692
rect 411 590 445 624
rect 411 522 445 556
rect 411 454 445 488
rect 411 386 445 420
rect 411 318 445 352
rect 411 250 445 284
rect 411 182 445 216
rect 411 114 445 148
rect 537 1066 571 1100
rect 537 998 571 1032
rect 537 930 571 964
rect 537 862 571 896
rect 537 794 571 828
rect 537 726 571 760
rect 537 658 571 692
rect 537 590 571 624
rect 537 522 571 556
rect 537 454 571 488
rect 537 386 571 420
rect 537 318 571 352
rect 537 250 571 284
rect 537 182 571 216
rect 537 114 571 148
rect 663 1066 697 1100
rect 663 998 697 1032
rect 663 930 697 964
rect 663 862 697 896
rect 663 794 697 828
rect 663 726 697 760
rect 663 658 697 692
rect 663 590 697 624
rect 663 522 697 556
rect 663 454 697 488
rect 663 386 697 420
rect 663 318 697 352
rect 663 250 697 284
rect 663 182 697 216
rect 663 114 697 148
<< nsubdiff >>
rect 36 1066 94 1112
rect 36 1032 48 1066
rect 82 1032 94 1066
rect 36 998 94 1032
rect 36 964 48 998
rect 82 964 94 998
rect 36 930 94 964
rect 36 896 48 930
rect 82 896 94 930
rect 36 862 94 896
rect 36 828 48 862
rect 82 828 94 862
rect 36 794 94 828
rect 36 760 48 794
rect 82 760 94 794
rect 36 726 94 760
rect 36 692 48 726
rect 82 692 94 726
rect 36 658 94 692
rect 36 624 48 658
rect 82 624 94 658
rect 36 590 94 624
rect 36 556 48 590
rect 82 556 94 590
rect 36 522 94 556
rect 36 488 48 522
rect 82 488 94 522
rect 36 454 94 488
rect 36 420 48 454
rect 82 420 94 454
rect 36 386 94 420
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 762 1066 820 1112
rect 762 1032 774 1066
rect 808 1032 820 1066
rect 762 998 820 1032
rect 762 964 774 998
rect 808 964 820 998
rect 762 930 820 964
rect 762 896 774 930
rect 808 896 820 930
rect 762 862 820 896
rect 762 828 774 862
rect 808 828 820 862
rect 762 794 820 828
rect 762 760 774 794
rect 808 760 820 794
rect 762 726 820 760
rect 762 692 774 726
rect 808 692 820 726
rect 762 658 820 692
rect 762 624 774 658
rect 808 624 820 658
rect 762 590 820 624
rect 762 556 774 590
rect 808 556 820 590
rect 762 522 820 556
rect 762 488 774 522
rect 808 488 820 522
rect 762 454 820 488
rect 762 420 774 454
rect 808 420 820 454
rect 762 386 820 420
rect 762 352 774 386
rect 808 352 820 386
rect 762 318 820 352
rect 762 284 774 318
rect 808 284 820 318
rect 762 250 820 284
rect 762 216 774 250
rect 808 216 820 250
rect 762 182 820 216
rect 762 148 774 182
rect 808 148 820 182
rect 762 102 820 148
<< nsubdiffcont >>
rect 48 1032 82 1066
rect 48 964 82 998
rect 48 896 82 930
rect 48 828 82 862
rect 48 760 82 794
rect 48 692 82 726
rect 48 624 82 658
rect 48 556 82 590
rect 48 488 82 522
rect 48 420 82 454
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 774 1032 808 1066
rect 774 964 808 998
rect 774 896 808 930
rect 774 828 808 862
rect 774 760 808 794
rect 774 692 808 726
rect 774 624 808 658
rect 774 556 808 590
rect 774 488 808 522
rect 774 420 808 454
rect 774 352 808 386
rect 774 284 808 318
rect 774 216 808 250
rect 774 148 808 182
<< poly >>
rect 191 1194 665 1214
rect 191 1160 207 1194
rect 241 1160 275 1194
rect 309 1160 343 1194
rect 377 1160 411 1194
rect 445 1160 479 1194
rect 513 1160 547 1194
rect 581 1160 615 1194
rect 649 1160 665 1194
rect 191 1144 665 1160
rect 204 1112 274 1144
rect 330 1112 400 1144
rect 456 1112 526 1144
rect 582 1112 652 1144
rect 204 70 274 102
rect 330 70 400 102
rect 456 70 526 102
rect 582 70 652 102
rect 191 54 665 70
rect 191 20 207 54
rect 241 20 275 54
rect 309 20 343 54
rect 377 20 411 54
rect 445 20 479 54
rect 513 20 547 54
rect 581 20 615 54
rect 649 20 665 54
rect 191 0 665 20
<< polycont >>
rect 207 1160 241 1194
rect 275 1160 309 1194
rect 343 1160 377 1194
rect 411 1160 445 1194
rect 479 1160 513 1194
rect 547 1160 581 1194
rect 615 1160 649 1194
rect 207 20 241 54
rect 275 20 309 54
rect 343 20 377 54
rect 411 20 445 54
rect 479 20 513 54
rect 547 20 581 54
rect 615 20 649 54
<< locali >>
rect 191 1160 195 1194
rect 241 1160 267 1194
rect 309 1160 339 1194
rect 377 1160 411 1194
rect 445 1160 479 1194
rect 517 1160 547 1194
rect 589 1160 615 1194
rect 661 1160 665 1194
rect 159 1100 193 1116
rect 48 1020 82 1032
rect 48 948 82 964
rect 48 876 82 896
rect 48 804 82 828
rect 48 732 82 760
rect 48 660 82 692
rect 48 590 82 624
rect 48 522 82 554
rect 48 454 82 482
rect 48 386 82 410
rect 48 318 82 338
rect 48 250 82 266
rect 48 182 82 194
rect 159 1032 193 1058
rect 159 964 193 986
rect 159 896 193 914
rect 159 828 193 842
rect 159 760 193 770
rect 159 692 193 698
rect 159 624 193 626
rect 159 588 193 590
rect 159 516 193 522
rect 159 444 193 454
rect 159 372 193 386
rect 159 300 193 318
rect 159 228 193 250
rect 159 156 193 182
rect 159 98 193 114
rect 285 1100 319 1116
rect 285 1032 319 1058
rect 285 964 319 986
rect 285 896 319 914
rect 285 828 319 842
rect 285 760 319 770
rect 285 692 319 698
rect 285 624 319 626
rect 285 588 319 590
rect 285 516 319 522
rect 285 444 319 454
rect 285 372 319 386
rect 285 300 319 318
rect 285 228 319 250
rect 285 156 319 182
rect 285 98 319 114
rect 411 1100 445 1116
rect 411 1032 445 1058
rect 411 964 445 986
rect 411 896 445 914
rect 411 828 445 842
rect 411 760 445 770
rect 411 692 445 698
rect 411 624 445 626
rect 411 588 445 590
rect 411 516 445 522
rect 411 444 445 454
rect 411 372 445 386
rect 411 300 445 318
rect 411 228 445 250
rect 411 156 445 182
rect 411 98 445 114
rect 537 1100 571 1116
rect 537 1032 571 1058
rect 537 964 571 986
rect 537 896 571 914
rect 537 828 571 842
rect 537 760 571 770
rect 537 692 571 698
rect 537 624 571 626
rect 537 588 571 590
rect 537 516 571 522
rect 537 444 571 454
rect 537 372 571 386
rect 537 300 571 318
rect 537 228 571 250
rect 537 156 571 182
rect 537 98 571 114
rect 663 1100 697 1116
rect 663 1032 697 1058
rect 663 964 697 986
rect 663 896 697 914
rect 663 828 697 842
rect 663 760 697 770
rect 663 692 697 698
rect 663 624 697 626
rect 663 588 697 590
rect 663 516 697 522
rect 663 444 697 454
rect 663 372 697 386
rect 663 300 697 318
rect 663 228 697 250
rect 663 156 697 182
rect 774 1020 808 1032
rect 774 948 808 964
rect 774 876 808 896
rect 774 804 808 828
rect 774 732 808 760
rect 774 660 808 692
rect 774 590 808 624
rect 774 522 808 554
rect 774 454 808 482
rect 774 386 808 410
rect 774 318 808 338
rect 774 250 808 266
rect 774 182 808 194
rect 663 98 697 114
rect 191 20 195 54
rect 241 20 267 54
rect 309 20 339 54
rect 377 20 411 54
rect 445 20 479 54
rect 517 20 547 54
rect 589 20 615 54
rect 661 20 665 54
<< viali >>
rect 195 1160 207 1194
rect 207 1160 229 1194
rect 267 1160 275 1194
rect 275 1160 301 1194
rect 339 1160 343 1194
rect 343 1160 373 1194
rect 411 1160 445 1194
rect 483 1160 513 1194
rect 513 1160 517 1194
rect 555 1160 581 1194
rect 581 1160 589 1194
rect 627 1160 649 1194
rect 649 1160 661 1194
rect 48 1066 82 1092
rect 48 1058 82 1066
rect 48 998 82 1020
rect 48 986 82 998
rect 48 930 82 948
rect 48 914 82 930
rect 48 862 82 876
rect 48 842 82 862
rect 48 794 82 804
rect 48 770 82 794
rect 48 726 82 732
rect 48 698 82 726
rect 48 658 82 660
rect 48 626 82 658
rect 48 556 82 588
rect 48 554 82 556
rect 48 488 82 516
rect 48 482 82 488
rect 48 420 82 444
rect 48 410 82 420
rect 48 352 82 372
rect 48 338 82 352
rect 48 284 82 300
rect 48 266 82 284
rect 48 216 82 228
rect 48 194 82 216
rect 48 148 82 156
rect 48 122 82 148
rect 159 1066 193 1092
rect 159 1058 193 1066
rect 159 998 193 1020
rect 159 986 193 998
rect 159 930 193 948
rect 159 914 193 930
rect 159 862 193 876
rect 159 842 193 862
rect 159 794 193 804
rect 159 770 193 794
rect 159 726 193 732
rect 159 698 193 726
rect 159 658 193 660
rect 159 626 193 658
rect 159 556 193 588
rect 159 554 193 556
rect 159 488 193 516
rect 159 482 193 488
rect 159 420 193 444
rect 159 410 193 420
rect 159 352 193 372
rect 159 338 193 352
rect 159 284 193 300
rect 159 266 193 284
rect 159 216 193 228
rect 159 194 193 216
rect 159 148 193 156
rect 159 122 193 148
rect 285 1066 319 1092
rect 285 1058 319 1066
rect 285 998 319 1020
rect 285 986 319 998
rect 285 930 319 948
rect 285 914 319 930
rect 285 862 319 876
rect 285 842 319 862
rect 285 794 319 804
rect 285 770 319 794
rect 285 726 319 732
rect 285 698 319 726
rect 285 658 319 660
rect 285 626 319 658
rect 285 556 319 588
rect 285 554 319 556
rect 285 488 319 516
rect 285 482 319 488
rect 285 420 319 444
rect 285 410 319 420
rect 285 352 319 372
rect 285 338 319 352
rect 285 284 319 300
rect 285 266 319 284
rect 285 216 319 228
rect 285 194 319 216
rect 285 148 319 156
rect 285 122 319 148
rect 411 1066 445 1092
rect 411 1058 445 1066
rect 411 998 445 1020
rect 411 986 445 998
rect 411 930 445 948
rect 411 914 445 930
rect 411 862 445 876
rect 411 842 445 862
rect 411 794 445 804
rect 411 770 445 794
rect 411 726 445 732
rect 411 698 445 726
rect 411 658 445 660
rect 411 626 445 658
rect 411 556 445 588
rect 411 554 445 556
rect 411 488 445 516
rect 411 482 445 488
rect 411 420 445 444
rect 411 410 445 420
rect 411 352 445 372
rect 411 338 445 352
rect 411 284 445 300
rect 411 266 445 284
rect 411 216 445 228
rect 411 194 445 216
rect 411 148 445 156
rect 411 122 445 148
rect 537 1066 571 1092
rect 537 1058 571 1066
rect 537 998 571 1020
rect 537 986 571 998
rect 537 930 571 948
rect 537 914 571 930
rect 537 862 571 876
rect 537 842 571 862
rect 537 794 571 804
rect 537 770 571 794
rect 537 726 571 732
rect 537 698 571 726
rect 537 658 571 660
rect 537 626 571 658
rect 537 556 571 588
rect 537 554 571 556
rect 537 488 571 516
rect 537 482 571 488
rect 537 420 571 444
rect 537 410 571 420
rect 537 352 571 372
rect 537 338 571 352
rect 537 284 571 300
rect 537 266 571 284
rect 537 216 571 228
rect 537 194 571 216
rect 537 148 571 156
rect 537 122 571 148
rect 663 1066 697 1092
rect 663 1058 697 1066
rect 663 998 697 1020
rect 663 986 697 998
rect 663 930 697 948
rect 663 914 697 930
rect 663 862 697 876
rect 663 842 697 862
rect 663 794 697 804
rect 663 770 697 794
rect 663 726 697 732
rect 663 698 697 726
rect 663 658 697 660
rect 663 626 697 658
rect 663 556 697 588
rect 663 554 697 556
rect 663 488 697 516
rect 663 482 697 488
rect 663 420 697 444
rect 663 410 697 420
rect 663 352 697 372
rect 663 338 697 352
rect 663 284 697 300
rect 663 266 697 284
rect 663 216 697 228
rect 663 194 697 216
rect 663 148 697 156
rect 663 122 697 148
rect 774 1066 808 1092
rect 774 1058 808 1066
rect 774 998 808 1020
rect 774 986 808 998
rect 774 930 808 948
rect 774 914 808 930
rect 774 862 808 876
rect 774 842 808 862
rect 774 794 808 804
rect 774 770 808 794
rect 774 726 808 732
rect 774 698 808 726
rect 774 658 808 660
rect 774 626 808 658
rect 774 556 808 588
rect 774 554 808 556
rect 774 488 808 516
rect 774 482 808 488
rect 774 420 808 444
rect 774 410 808 420
rect 774 352 808 372
rect 774 338 808 352
rect 774 284 808 300
rect 774 266 808 284
rect 774 216 808 228
rect 774 194 808 216
rect 774 148 808 156
rect 774 122 808 148
rect 195 20 207 54
rect 207 20 229 54
rect 267 20 275 54
rect 275 20 301 54
rect 339 20 343 54
rect 343 20 373 54
rect 411 20 445 54
rect 483 20 513 54
rect 513 20 517 54
rect 555 20 581 54
rect 581 20 589 54
rect 627 20 649 54
rect 649 20 661 54
<< metal1 >>
rect 183 1194 673 1214
rect 183 1160 195 1194
rect 229 1160 267 1194
rect 301 1160 339 1194
rect 373 1160 411 1194
rect 445 1160 483 1194
rect 517 1160 555 1194
rect 589 1160 627 1194
rect 661 1160 673 1194
rect 183 1148 673 1160
rect 36 1092 94 1104
rect 36 1058 48 1092
rect 82 1058 94 1092
rect 36 1020 94 1058
rect 36 986 48 1020
rect 82 986 94 1020
rect 36 948 94 986
rect 36 914 48 948
rect 82 914 94 948
rect 36 876 94 914
rect 36 842 48 876
rect 82 842 94 876
rect 36 804 94 842
rect 36 770 48 804
rect 82 770 94 804
rect 36 732 94 770
rect 36 698 48 732
rect 82 698 94 732
rect 36 660 94 698
rect 36 626 48 660
rect 82 626 94 660
rect 36 588 94 626
rect 36 554 48 588
rect 82 554 94 588
rect 36 516 94 554
rect 36 482 48 516
rect 82 482 94 516
rect 36 444 94 482
rect 36 410 48 444
rect 82 410 94 444
rect 36 372 94 410
rect 36 338 48 372
rect 82 338 94 372
rect 36 300 94 338
rect 36 266 48 300
rect 82 266 94 300
rect 36 228 94 266
rect 36 194 48 228
rect 82 194 94 228
rect 36 156 94 194
rect 36 122 48 156
rect 82 122 94 156
rect 36 110 94 122
rect 150 1092 202 1104
rect 150 1058 159 1092
rect 193 1058 202 1092
rect 150 1020 202 1058
rect 150 986 159 1020
rect 193 986 202 1020
rect 150 948 202 986
rect 150 914 159 948
rect 193 914 202 948
rect 150 876 202 914
rect 150 842 159 876
rect 193 842 202 876
rect 150 804 202 842
rect 150 770 159 804
rect 193 770 202 804
rect 150 732 202 770
rect 150 698 159 732
rect 193 698 202 732
rect 150 660 202 698
rect 150 626 159 660
rect 193 626 202 660
rect 150 588 202 626
rect 150 554 159 588
rect 193 554 202 588
rect 150 552 202 554
rect 150 488 159 500
rect 193 488 202 500
rect 150 424 159 436
rect 193 424 202 436
rect 150 360 159 372
rect 193 360 202 372
rect 150 300 202 308
rect 150 296 159 300
rect 193 296 202 300
rect 150 232 202 244
rect 150 168 202 180
rect 150 110 202 116
rect 276 1098 328 1104
rect 276 1034 328 1046
rect 276 970 328 982
rect 276 914 285 918
rect 319 914 328 918
rect 276 906 328 914
rect 276 842 285 854
rect 319 842 328 854
rect 276 778 285 790
rect 319 778 328 790
rect 276 714 285 726
rect 319 714 328 726
rect 276 660 328 662
rect 276 626 285 660
rect 319 626 328 660
rect 276 588 328 626
rect 276 554 285 588
rect 319 554 328 588
rect 276 516 328 554
rect 276 482 285 516
rect 319 482 328 516
rect 276 444 328 482
rect 276 410 285 444
rect 319 410 328 444
rect 276 372 328 410
rect 276 338 285 372
rect 319 338 328 372
rect 276 300 328 338
rect 276 266 285 300
rect 319 266 328 300
rect 276 228 328 266
rect 276 194 285 228
rect 319 194 328 228
rect 276 156 328 194
rect 276 122 285 156
rect 319 122 328 156
rect 276 110 328 122
rect 402 1092 454 1104
rect 402 1058 411 1092
rect 445 1058 454 1092
rect 402 1020 454 1058
rect 402 986 411 1020
rect 445 986 454 1020
rect 402 948 454 986
rect 402 914 411 948
rect 445 914 454 948
rect 402 876 454 914
rect 402 842 411 876
rect 445 842 454 876
rect 402 804 454 842
rect 402 770 411 804
rect 445 770 454 804
rect 402 732 454 770
rect 402 698 411 732
rect 445 698 454 732
rect 402 660 454 698
rect 402 626 411 660
rect 445 626 454 660
rect 402 588 454 626
rect 402 554 411 588
rect 445 554 454 588
rect 402 552 454 554
rect 402 488 411 500
rect 445 488 454 500
rect 402 424 411 436
rect 445 424 454 436
rect 402 360 411 372
rect 445 360 454 372
rect 402 300 454 308
rect 402 296 411 300
rect 445 296 454 300
rect 402 232 454 244
rect 402 168 454 180
rect 402 110 454 116
rect 528 1098 580 1104
rect 528 1034 580 1046
rect 528 970 580 982
rect 528 914 537 918
rect 571 914 580 918
rect 528 906 580 914
rect 528 842 537 854
rect 571 842 580 854
rect 528 778 537 790
rect 571 778 580 790
rect 528 714 537 726
rect 571 714 580 726
rect 528 660 580 662
rect 528 626 537 660
rect 571 626 580 660
rect 528 588 580 626
rect 528 554 537 588
rect 571 554 580 588
rect 528 516 580 554
rect 528 482 537 516
rect 571 482 580 516
rect 528 444 580 482
rect 528 410 537 444
rect 571 410 580 444
rect 528 372 580 410
rect 528 338 537 372
rect 571 338 580 372
rect 528 300 580 338
rect 528 266 537 300
rect 571 266 580 300
rect 528 228 580 266
rect 528 194 537 228
rect 571 194 580 228
rect 528 156 580 194
rect 528 122 537 156
rect 571 122 580 156
rect 528 110 580 122
rect 654 1092 706 1104
rect 654 1058 663 1092
rect 697 1058 706 1092
rect 654 1020 706 1058
rect 654 986 663 1020
rect 697 986 706 1020
rect 654 948 706 986
rect 654 914 663 948
rect 697 914 706 948
rect 654 876 706 914
rect 654 842 663 876
rect 697 842 706 876
rect 654 804 706 842
rect 654 770 663 804
rect 697 770 706 804
rect 654 732 706 770
rect 654 698 663 732
rect 697 698 706 732
rect 654 660 706 698
rect 654 626 663 660
rect 697 626 706 660
rect 654 588 706 626
rect 654 554 663 588
rect 697 554 706 588
rect 654 552 706 554
rect 654 488 663 500
rect 697 488 706 500
rect 654 424 663 436
rect 697 424 706 436
rect 654 360 663 372
rect 697 360 706 372
rect 654 300 706 308
rect 654 296 663 300
rect 697 296 706 300
rect 654 232 706 244
rect 654 168 706 180
rect 654 110 706 116
rect 762 1092 820 1104
rect 762 1058 774 1092
rect 808 1058 820 1092
rect 762 1020 820 1058
rect 762 986 774 1020
rect 808 986 820 1020
rect 762 948 820 986
rect 762 914 774 948
rect 808 914 820 948
rect 762 876 820 914
rect 762 842 774 876
rect 808 842 820 876
rect 762 804 820 842
rect 762 770 774 804
rect 808 770 820 804
rect 762 732 820 770
rect 762 698 774 732
rect 808 698 820 732
rect 762 660 820 698
rect 762 626 774 660
rect 808 626 820 660
rect 762 588 820 626
rect 762 554 774 588
rect 808 554 820 588
rect 762 516 820 554
rect 762 482 774 516
rect 808 482 820 516
rect 762 444 820 482
rect 762 410 774 444
rect 808 410 820 444
rect 762 372 820 410
rect 762 338 774 372
rect 808 338 820 372
rect 762 300 820 338
rect 762 266 774 300
rect 808 266 820 300
rect 762 228 820 266
rect 762 194 774 228
rect 808 194 820 228
rect 762 156 820 194
rect 762 122 774 156
rect 808 122 820 156
rect 762 110 820 122
rect 183 54 673 66
rect 183 20 195 54
rect 229 20 267 54
rect 301 20 339 54
rect 373 20 411 54
rect 445 20 483 54
rect 517 20 555 54
rect 589 20 627 54
rect 661 20 673 54
rect 183 0 673 20
<< via1 >>
rect 150 516 202 552
rect 150 500 159 516
rect 159 500 193 516
rect 193 500 202 516
rect 150 482 159 488
rect 159 482 193 488
rect 193 482 202 488
rect 150 444 202 482
rect 150 436 159 444
rect 159 436 193 444
rect 193 436 202 444
rect 150 410 159 424
rect 159 410 193 424
rect 193 410 202 424
rect 150 372 202 410
rect 150 338 159 360
rect 159 338 193 360
rect 193 338 202 360
rect 150 308 202 338
rect 150 266 159 296
rect 159 266 193 296
rect 193 266 202 296
rect 150 244 202 266
rect 150 228 202 232
rect 150 194 159 228
rect 159 194 193 228
rect 193 194 202 228
rect 150 180 202 194
rect 150 156 202 168
rect 150 122 159 156
rect 159 122 193 156
rect 193 122 202 156
rect 150 116 202 122
rect 276 1092 328 1098
rect 276 1058 285 1092
rect 285 1058 319 1092
rect 319 1058 328 1092
rect 276 1046 328 1058
rect 276 1020 328 1034
rect 276 986 285 1020
rect 285 986 319 1020
rect 319 986 328 1020
rect 276 982 328 986
rect 276 948 328 970
rect 276 918 285 948
rect 285 918 319 948
rect 319 918 328 948
rect 276 876 328 906
rect 276 854 285 876
rect 285 854 319 876
rect 319 854 328 876
rect 276 804 328 842
rect 276 790 285 804
rect 285 790 319 804
rect 319 790 328 804
rect 276 770 285 778
rect 285 770 319 778
rect 319 770 328 778
rect 276 732 328 770
rect 276 726 285 732
rect 285 726 319 732
rect 319 726 328 732
rect 276 698 285 714
rect 285 698 319 714
rect 319 698 328 714
rect 276 662 328 698
rect 402 516 454 552
rect 402 500 411 516
rect 411 500 445 516
rect 445 500 454 516
rect 402 482 411 488
rect 411 482 445 488
rect 445 482 454 488
rect 402 444 454 482
rect 402 436 411 444
rect 411 436 445 444
rect 445 436 454 444
rect 402 410 411 424
rect 411 410 445 424
rect 445 410 454 424
rect 402 372 454 410
rect 402 338 411 360
rect 411 338 445 360
rect 445 338 454 360
rect 402 308 454 338
rect 402 266 411 296
rect 411 266 445 296
rect 445 266 454 296
rect 402 244 454 266
rect 402 228 454 232
rect 402 194 411 228
rect 411 194 445 228
rect 445 194 454 228
rect 402 180 454 194
rect 402 156 454 168
rect 402 122 411 156
rect 411 122 445 156
rect 445 122 454 156
rect 402 116 454 122
rect 528 1092 580 1098
rect 528 1058 537 1092
rect 537 1058 571 1092
rect 571 1058 580 1092
rect 528 1046 580 1058
rect 528 1020 580 1034
rect 528 986 537 1020
rect 537 986 571 1020
rect 571 986 580 1020
rect 528 982 580 986
rect 528 948 580 970
rect 528 918 537 948
rect 537 918 571 948
rect 571 918 580 948
rect 528 876 580 906
rect 528 854 537 876
rect 537 854 571 876
rect 571 854 580 876
rect 528 804 580 842
rect 528 790 537 804
rect 537 790 571 804
rect 571 790 580 804
rect 528 770 537 778
rect 537 770 571 778
rect 571 770 580 778
rect 528 732 580 770
rect 528 726 537 732
rect 537 726 571 732
rect 571 726 580 732
rect 528 698 537 714
rect 537 698 571 714
rect 571 698 580 714
rect 528 662 580 698
rect 654 516 706 552
rect 654 500 663 516
rect 663 500 697 516
rect 697 500 706 516
rect 654 482 663 488
rect 663 482 697 488
rect 697 482 706 488
rect 654 444 706 482
rect 654 436 663 444
rect 663 436 697 444
rect 697 436 706 444
rect 654 410 663 424
rect 663 410 697 424
rect 697 410 706 424
rect 654 372 706 410
rect 654 338 663 360
rect 663 338 697 360
rect 697 338 706 360
rect 654 308 706 338
rect 654 266 663 296
rect 663 266 697 296
rect 697 266 706 296
rect 654 244 706 266
rect 654 228 706 232
rect 654 194 663 228
rect 663 194 697 228
rect 697 194 706 228
rect 654 180 706 194
rect 654 156 706 168
rect 654 122 663 156
rect 663 122 697 156
rect 697 122 706 156
rect 654 116 706 122
<< metal2 >>
rect 10 1098 846 1104
rect 10 1046 276 1098
rect 328 1046 528 1098
rect 580 1046 846 1098
rect 10 1034 846 1046
rect 10 982 276 1034
rect 328 982 528 1034
rect 580 982 846 1034
rect 10 970 846 982
rect 10 918 276 970
rect 328 918 528 970
rect 580 918 846 970
rect 10 906 846 918
rect 10 854 276 906
rect 328 854 528 906
rect 580 854 846 906
rect 10 842 846 854
rect 10 790 276 842
rect 328 790 528 842
rect 580 790 846 842
rect 10 778 846 790
rect 10 726 276 778
rect 328 726 528 778
rect 580 726 846 778
rect 10 714 846 726
rect 10 662 276 714
rect 328 662 528 714
rect 580 662 846 714
rect 10 632 846 662
rect 10 552 846 582
rect 10 500 150 552
rect 202 500 402 552
rect 454 500 654 552
rect 706 500 846 552
rect 10 488 846 500
rect 10 436 150 488
rect 202 436 402 488
rect 454 436 654 488
rect 706 436 846 488
rect 10 424 846 436
rect 10 372 150 424
rect 202 372 402 424
rect 454 372 654 424
rect 706 372 846 424
rect 10 360 846 372
rect 10 308 150 360
rect 202 308 402 360
rect 454 308 654 360
rect 706 308 846 360
rect 10 296 846 308
rect 10 244 150 296
rect 202 244 402 296
rect 454 244 654 296
rect 706 244 846 296
rect 10 232 846 244
rect 10 180 150 232
rect 202 180 402 232
rect 454 180 654 232
rect 706 180 846 232
rect 10 168 846 180
rect 10 116 150 168
rect 202 116 402 168
rect 454 116 654 168
rect 706 116 846 168
rect 10 110 846 116
<< labels >>
flabel metal2 s 15 798 34 868 0 FreeSans 400 90 0 0 DRAIN
port 2 nsew
flabel metal2 s 14 317 35 381 0 FreeSans 400 90 0 0 SOURCE
port 3 nsew
flabel metal1 s 60 730 60 730 7 FreeSans 400 90 0 0 BULK
flabel metal1 s 790 730 790 730 7 FreeSans 400 90 0 0 BULK
flabel metal1 s 183 1148 673 1214 0 FreeSans 300 0 0 0 GATE
port 4 nsew
flabel metal1 s 183 0 673 66 0 FreeSans 300 0 0 0 GATE
port 4 nsew
<< properties >>
string GDS_END 10001302
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9979334
<< end >>
