magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< metal3 >>
rect 120 3272 4900 3276
rect 120 3208 126 3272
rect 190 3208 208 3272
rect 272 3208 290 3272
rect 354 3208 372 3272
rect 436 3208 454 3272
rect 518 3208 536 3272
rect 600 3208 618 3272
rect 682 3208 699 3272
rect 763 3208 780 3272
rect 844 3208 861 3272
rect 925 3208 942 3272
rect 1006 3208 1023 3272
rect 1087 3208 1104 3272
rect 1168 3208 1185 3272
rect 1249 3208 1266 3272
rect 1330 3208 1347 3272
rect 1411 3208 1428 3272
rect 1492 3208 1509 3272
rect 1573 3208 1590 3272
rect 1654 3208 1671 3272
rect 1735 3208 1752 3272
rect 1816 3208 1833 3272
rect 1897 3208 1914 3272
rect 1978 3208 1995 3272
rect 2059 3208 2076 3272
rect 2140 3208 2157 3272
rect 2221 3208 2238 3272
rect 2302 3208 2319 3272
rect 2383 3208 2400 3272
rect 2464 3208 2481 3272
rect 2545 3208 2562 3272
rect 2626 3208 2643 3272
rect 2707 3208 2724 3272
rect 2788 3208 2805 3272
rect 2869 3208 2886 3272
rect 2950 3208 2967 3272
rect 3031 3208 3048 3272
rect 3112 3208 3129 3272
rect 3193 3208 3210 3272
rect 3274 3208 3291 3272
rect 3355 3208 3372 3272
rect 3436 3208 3453 3272
rect 3517 3208 3534 3272
rect 3598 3208 3615 3272
rect 3679 3208 3696 3272
rect 3760 3208 3777 3272
rect 3841 3208 3858 3272
rect 3922 3208 3939 3272
rect 4003 3208 4020 3272
rect 4084 3208 4101 3272
rect 4165 3208 4182 3272
rect 4246 3208 4263 3272
rect 4327 3208 4344 3272
rect 4408 3208 4425 3272
rect 4489 3208 4506 3272
rect 4570 3208 4587 3272
rect 4651 3208 4668 3272
rect 4732 3208 4749 3272
rect 4813 3208 4830 3272
rect 4894 3208 4900 3272
rect 120 3184 4900 3208
rect 120 3120 126 3184
rect 190 3120 208 3184
rect 272 3120 290 3184
rect 354 3120 372 3184
rect 436 3120 454 3184
rect 518 3120 536 3184
rect 600 3120 618 3184
rect 682 3120 699 3184
rect 763 3120 780 3184
rect 844 3120 861 3184
rect 925 3120 942 3184
rect 1006 3120 1023 3184
rect 1087 3120 1104 3184
rect 1168 3120 1185 3184
rect 1249 3120 1266 3184
rect 1330 3120 1347 3184
rect 1411 3120 1428 3184
rect 1492 3120 1509 3184
rect 1573 3120 1590 3184
rect 1654 3120 1671 3184
rect 1735 3120 1752 3184
rect 1816 3120 1833 3184
rect 1897 3120 1914 3184
rect 1978 3120 1995 3184
rect 2059 3120 2076 3184
rect 2140 3120 2157 3184
rect 2221 3120 2238 3184
rect 2302 3120 2319 3184
rect 2383 3120 2400 3184
rect 2464 3120 2481 3184
rect 2545 3120 2562 3184
rect 2626 3120 2643 3184
rect 2707 3120 2724 3184
rect 2788 3120 2805 3184
rect 2869 3120 2886 3184
rect 2950 3120 2967 3184
rect 3031 3120 3048 3184
rect 3112 3120 3129 3184
rect 3193 3120 3210 3184
rect 3274 3120 3291 3184
rect 3355 3120 3372 3184
rect 3436 3120 3453 3184
rect 3517 3120 3534 3184
rect 3598 3120 3615 3184
rect 3679 3120 3696 3184
rect 3760 3120 3777 3184
rect 3841 3120 3858 3184
rect 3922 3120 3939 3184
rect 4003 3120 4020 3184
rect 4084 3120 4101 3184
rect 4165 3120 4182 3184
rect 4246 3120 4263 3184
rect 4327 3120 4344 3184
rect 4408 3120 4425 3184
rect 4489 3120 4506 3184
rect 4570 3120 4587 3184
rect 4651 3120 4668 3184
rect 4732 3120 4749 3184
rect 4813 3120 4830 3184
rect 4894 3120 4900 3184
rect 120 3096 4900 3120
rect 120 3032 126 3096
rect 190 3032 208 3096
rect 272 3032 290 3096
rect 354 3032 372 3096
rect 436 3032 454 3096
rect 518 3032 536 3096
rect 600 3032 618 3096
rect 682 3032 699 3096
rect 763 3032 780 3096
rect 844 3032 861 3096
rect 925 3032 942 3096
rect 1006 3032 1023 3096
rect 1087 3032 1104 3096
rect 1168 3032 1185 3096
rect 1249 3032 1266 3096
rect 1330 3032 1347 3096
rect 1411 3032 1428 3096
rect 1492 3032 1509 3096
rect 1573 3032 1590 3096
rect 1654 3032 1671 3096
rect 1735 3032 1752 3096
rect 1816 3032 1833 3096
rect 1897 3032 1914 3096
rect 1978 3032 1995 3096
rect 2059 3032 2076 3096
rect 2140 3032 2157 3096
rect 2221 3032 2238 3096
rect 2302 3032 2319 3096
rect 2383 3032 2400 3096
rect 2464 3032 2481 3096
rect 2545 3032 2562 3096
rect 2626 3032 2643 3096
rect 2707 3032 2724 3096
rect 2788 3032 2805 3096
rect 2869 3032 2886 3096
rect 2950 3032 2967 3096
rect 3031 3032 3048 3096
rect 3112 3032 3129 3096
rect 3193 3032 3210 3096
rect 3274 3032 3291 3096
rect 3355 3032 3372 3096
rect 3436 3032 3453 3096
rect 3517 3032 3534 3096
rect 3598 3032 3615 3096
rect 3679 3032 3696 3096
rect 3760 3032 3777 3096
rect 3841 3032 3858 3096
rect 3922 3032 3939 3096
rect 4003 3032 4020 3096
rect 4084 3032 4101 3096
rect 4165 3032 4182 3096
rect 4246 3032 4263 3096
rect 4327 3032 4344 3096
rect 4408 3032 4425 3096
rect 4489 3032 4506 3096
rect 4570 3032 4587 3096
rect 4651 3032 4668 3096
rect 4732 3032 4749 3096
rect 4813 3032 4830 3096
rect 4894 3032 4900 3096
rect 120 3008 4900 3032
rect 120 2944 126 3008
rect 190 2944 208 3008
rect 272 2944 290 3008
rect 354 2944 372 3008
rect 436 2944 454 3008
rect 518 2944 536 3008
rect 600 2944 618 3008
rect 682 2944 699 3008
rect 763 2944 780 3008
rect 844 2944 861 3008
rect 925 2944 942 3008
rect 1006 2944 1023 3008
rect 1087 2944 1104 3008
rect 1168 2944 1185 3008
rect 1249 2944 1266 3008
rect 1330 2944 1347 3008
rect 1411 2944 1428 3008
rect 1492 2944 1509 3008
rect 1573 2944 1590 3008
rect 1654 2944 1671 3008
rect 1735 2944 1752 3008
rect 1816 2944 1833 3008
rect 1897 2944 1914 3008
rect 1978 2944 1995 3008
rect 2059 2944 2076 3008
rect 2140 2944 2157 3008
rect 2221 2944 2238 3008
rect 2302 2944 2319 3008
rect 2383 2944 2400 3008
rect 2464 2944 2481 3008
rect 2545 2944 2562 3008
rect 2626 2944 2643 3008
rect 2707 2944 2724 3008
rect 2788 2944 2805 3008
rect 2869 2944 2886 3008
rect 2950 2944 2967 3008
rect 3031 2944 3048 3008
rect 3112 2944 3129 3008
rect 3193 2944 3210 3008
rect 3274 2944 3291 3008
rect 3355 2944 3372 3008
rect 3436 2944 3453 3008
rect 3517 2944 3534 3008
rect 3598 2944 3615 3008
rect 3679 2944 3696 3008
rect 3760 2944 3777 3008
rect 3841 2944 3858 3008
rect 3922 2944 3939 3008
rect 4003 2944 4020 3008
rect 4084 2944 4101 3008
rect 4165 2944 4182 3008
rect 4246 2944 4263 3008
rect 4327 2944 4344 3008
rect 4408 2944 4425 3008
rect 4489 2944 4506 3008
rect 4570 2944 4587 3008
rect 4651 2944 4668 3008
rect 4732 2944 4749 3008
rect 4813 2944 4830 3008
rect 4894 2944 4900 3008
rect 120 2920 4900 2944
rect 120 2856 126 2920
rect 190 2856 208 2920
rect 272 2856 290 2920
rect 354 2856 372 2920
rect 436 2856 454 2920
rect 518 2856 536 2920
rect 600 2856 618 2920
rect 682 2856 699 2920
rect 763 2856 780 2920
rect 844 2856 861 2920
rect 925 2856 942 2920
rect 1006 2856 1023 2920
rect 1087 2856 1104 2920
rect 1168 2856 1185 2920
rect 1249 2856 1266 2920
rect 1330 2856 1347 2920
rect 1411 2856 1428 2920
rect 1492 2856 1509 2920
rect 1573 2856 1590 2920
rect 1654 2856 1671 2920
rect 1735 2856 1752 2920
rect 1816 2856 1833 2920
rect 1897 2856 1914 2920
rect 1978 2856 1995 2920
rect 2059 2856 2076 2920
rect 2140 2856 2157 2920
rect 2221 2856 2238 2920
rect 2302 2856 2319 2920
rect 2383 2856 2400 2920
rect 2464 2856 2481 2920
rect 2545 2856 2562 2920
rect 2626 2856 2643 2920
rect 2707 2856 2724 2920
rect 2788 2856 2805 2920
rect 2869 2856 2886 2920
rect 2950 2856 2967 2920
rect 3031 2856 3048 2920
rect 3112 2856 3129 2920
rect 3193 2856 3210 2920
rect 3274 2856 3291 2920
rect 3355 2856 3372 2920
rect 3436 2856 3453 2920
rect 3517 2856 3534 2920
rect 3598 2856 3615 2920
rect 3679 2856 3696 2920
rect 3760 2856 3777 2920
rect 3841 2856 3858 2920
rect 3922 2856 3939 2920
rect 4003 2856 4020 2920
rect 4084 2856 4101 2920
rect 4165 2856 4182 2920
rect 4246 2856 4263 2920
rect 4327 2856 4344 2920
rect 4408 2856 4425 2920
rect 4489 2856 4506 2920
rect 4570 2856 4587 2920
rect 4651 2856 4668 2920
rect 4732 2856 4749 2920
rect 4813 2856 4830 2920
rect 4894 2856 4900 2920
rect 120 2832 4900 2856
rect 120 2768 126 2832
rect 190 2768 208 2832
rect 272 2768 290 2832
rect 354 2768 372 2832
rect 436 2768 454 2832
rect 518 2768 536 2832
rect 600 2768 618 2832
rect 682 2768 699 2832
rect 763 2768 780 2832
rect 844 2768 861 2832
rect 925 2768 942 2832
rect 1006 2768 1023 2832
rect 1087 2768 1104 2832
rect 1168 2768 1185 2832
rect 1249 2768 1266 2832
rect 1330 2768 1347 2832
rect 1411 2768 1428 2832
rect 1492 2768 1509 2832
rect 1573 2768 1590 2832
rect 1654 2768 1671 2832
rect 1735 2768 1752 2832
rect 1816 2768 1833 2832
rect 1897 2768 1914 2832
rect 1978 2768 1995 2832
rect 2059 2768 2076 2832
rect 2140 2768 2157 2832
rect 2221 2768 2238 2832
rect 2302 2768 2319 2832
rect 2383 2768 2400 2832
rect 2464 2768 2481 2832
rect 2545 2768 2562 2832
rect 2626 2768 2643 2832
rect 2707 2768 2724 2832
rect 2788 2768 2805 2832
rect 2869 2768 2886 2832
rect 2950 2768 2967 2832
rect 3031 2768 3048 2832
rect 3112 2768 3129 2832
rect 3193 2768 3210 2832
rect 3274 2768 3291 2832
rect 3355 2768 3372 2832
rect 3436 2768 3453 2832
rect 3517 2768 3534 2832
rect 3598 2768 3615 2832
rect 3679 2768 3696 2832
rect 3760 2768 3777 2832
rect 3841 2768 3858 2832
rect 3922 2768 3939 2832
rect 4003 2768 4020 2832
rect 4084 2768 4101 2832
rect 4165 2768 4182 2832
rect 4246 2768 4263 2832
rect 4327 2768 4344 2832
rect 4408 2768 4425 2832
rect 4489 2768 4506 2832
rect 4570 2768 4587 2832
rect 4651 2768 4668 2832
rect 4732 2768 4749 2832
rect 4813 2768 4830 2832
rect 4894 2768 4900 2832
rect 120 2744 4900 2768
rect 120 2680 126 2744
rect 190 2680 208 2744
rect 272 2680 290 2744
rect 354 2680 372 2744
rect 436 2680 454 2744
rect 518 2680 536 2744
rect 600 2680 618 2744
rect 682 2680 699 2744
rect 763 2680 780 2744
rect 844 2680 861 2744
rect 925 2680 942 2744
rect 1006 2680 1023 2744
rect 1087 2680 1104 2744
rect 1168 2680 1185 2744
rect 1249 2680 1266 2744
rect 1330 2680 1347 2744
rect 1411 2680 1428 2744
rect 1492 2680 1509 2744
rect 1573 2680 1590 2744
rect 1654 2680 1671 2744
rect 1735 2680 1752 2744
rect 1816 2680 1833 2744
rect 1897 2680 1914 2744
rect 1978 2680 1995 2744
rect 2059 2680 2076 2744
rect 2140 2680 2157 2744
rect 2221 2680 2238 2744
rect 2302 2680 2319 2744
rect 2383 2680 2400 2744
rect 2464 2680 2481 2744
rect 2545 2680 2562 2744
rect 2626 2680 2643 2744
rect 2707 2680 2724 2744
rect 2788 2680 2805 2744
rect 2869 2680 2886 2744
rect 2950 2680 2967 2744
rect 3031 2680 3048 2744
rect 3112 2680 3129 2744
rect 3193 2680 3210 2744
rect 3274 2680 3291 2744
rect 3355 2680 3372 2744
rect 3436 2680 3453 2744
rect 3517 2680 3534 2744
rect 3598 2680 3615 2744
rect 3679 2680 3696 2744
rect 3760 2680 3777 2744
rect 3841 2680 3858 2744
rect 3922 2680 3939 2744
rect 4003 2680 4020 2744
rect 4084 2680 4101 2744
rect 4165 2680 4182 2744
rect 4246 2680 4263 2744
rect 4327 2680 4344 2744
rect 4408 2680 4425 2744
rect 4489 2680 4506 2744
rect 4570 2680 4587 2744
rect 4651 2680 4668 2744
rect 4732 2680 4749 2744
rect 4813 2680 4830 2744
rect 4894 2680 4900 2744
rect 120 2656 4900 2680
rect 120 2592 126 2656
rect 190 2592 208 2656
rect 272 2592 290 2656
rect 354 2592 372 2656
rect 436 2592 454 2656
rect 518 2592 536 2656
rect 600 2592 618 2656
rect 682 2592 699 2656
rect 763 2592 780 2656
rect 844 2592 861 2656
rect 925 2592 942 2656
rect 1006 2592 1023 2656
rect 1087 2592 1104 2656
rect 1168 2592 1185 2656
rect 1249 2592 1266 2656
rect 1330 2592 1347 2656
rect 1411 2592 1428 2656
rect 1492 2592 1509 2656
rect 1573 2592 1590 2656
rect 1654 2592 1671 2656
rect 1735 2592 1752 2656
rect 1816 2592 1833 2656
rect 1897 2592 1914 2656
rect 1978 2592 1995 2656
rect 2059 2592 2076 2656
rect 2140 2592 2157 2656
rect 2221 2592 2238 2656
rect 2302 2592 2319 2656
rect 2383 2592 2400 2656
rect 2464 2592 2481 2656
rect 2545 2592 2562 2656
rect 2626 2592 2643 2656
rect 2707 2592 2724 2656
rect 2788 2592 2805 2656
rect 2869 2592 2886 2656
rect 2950 2592 2967 2656
rect 3031 2592 3048 2656
rect 3112 2592 3129 2656
rect 3193 2592 3210 2656
rect 3274 2592 3291 2656
rect 3355 2592 3372 2656
rect 3436 2592 3453 2656
rect 3517 2592 3534 2656
rect 3598 2592 3615 2656
rect 3679 2592 3696 2656
rect 3760 2592 3777 2656
rect 3841 2592 3858 2656
rect 3922 2592 3939 2656
rect 4003 2592 4020 2656
rect 4084 2592 4101 2656
rect 4165 2592 4182 2656
rect 4246 2592 4263 2656
rect 4327 2592 4344 2656
rect 4408 2592 4425 2656
rect 4489 2592 4506 2656
rect 4570 2592 4587 2656
rect 4651 2592 4668 2656
rect 4732 2592 4749 2656
rect 4813 2592 4830 2656
rect 4894 2592 4900 2656
rect 120 2588 4900 2592
rect 10151 3272 14931 3276
rect 10151 3208 10157 3272
rect 10221 3208 10239 3272
rect 10303 3208 10321 3272
rect 10385 3208 10403 3272
rect 10467 3208 10485 3272
rect 10549 3208 10567 3272
rect 10631 3208 10649 3272
rect 10713 3208 10730 3272
rect 10794 3208 10811 3272
rect 10875 3208 10892 3272
rect 10956 3208 10973 3272
rect 11037 3208 11054 3272
rect 11118 3208 11135 3272
rect 11199 3208 11216 3272
rect 11280 3208 11297 3272
rect 11361 3208 11378 3272
rect 11442 3208 11459 3272
rect 11523 3208 11540 3272
rect 11604 3208 11621 3272
rect 11685 3208 11702 3272
rect 11766 3208 11783 3272
rect 11847 3208 11864 3272
rect 11928 3208 11945 3272
rect 12009 3208 12026 3272
rect 12090 3208 12107 3272
rect 12171 3208 12188 3272
rect 12252 3208 12269 3272
rect 12333 3208 12350 3272
rect 12414 3208 12431 3272
rect 12495 3208 12512 3272
rect 12576 3208 12593 3272
rect 12657 3208 12674 3272
rect 12738 3208 12755 3272
rect 12819 3208 12836 3272
rect 12900 3208 12917 3272
rect 12981 3208 12998 3272
rect 13062 3208 13079 3272
rect 13143 3208 13160 3272
rect 13224 3208 13241 3272
rect 13305 3208 13322 3272
rect 13386 3208 13403 3272
rect 13467 3208 13484 3272
rect 13548 3208 13565 3272
rect 13629 3208 13646 3272
rect 13710 3208 13727 3272
rect 13791 3208 13808 3272
rect 13872 3208 13889 3272
rect 13953 3208 13970 3272
rect 14034 3208 14051 3272
rect 14115 3208 14132 3272
rect 14196 3208 14213 3272
rect 14277 3208 14294 3272
rect 14358 3208 14375 3272
rect 14439 3208 14456 3272
rect 14520 3208 14537 3272
rect 14601 3208 14618 3272
rect 14682 3208 14699 3272
rect 14763 3208 14780 3272
rect 14844 3208 14861 3272
rect 14925 3208 14931 3272
rect 10151 3184 14931 3208
rect 10151 3120 10157 3184
rect 10221 3120 10239 3184
rect 10303 3120 10321 3184
rect 10385 3120 10403 3184
rect 10467 3120 10485 3184
rect 10549 3120 10567 3184
rect 10631 3120 10649 3184
rect 10713 3120 10730 3184
rect 10794 3120 10811 3184
rect 10875 3120 10892 3184
rect 10956 3120 10973 3184
rect 11037 3120 11054 3184
rect 11118 3120 11135 3184
rect 11199 3120 11216 3184
rect 11280 3120 11297 3184
rect 11361 3120 11378 3184
rect 11442 3120 11459 3184
rect 11523 3120 11540 3184
rect 11604 3120 11621 3184
rect 11685 3120 11702 3184
rect 11766 3120 11783 3184
rect 11847 3120 11864 3184
rect 11928 3120 11945 3184
rect 12009 3120 12026 3184
rect 12090 3120 12107 3184
rect 12171 3120 12188 3184
rect 12252 3120 12269 3184
rect 12333 3120 12350 3184
rect 12414 3120 12431 3184
rect 12495 3120 12512 3184
rect 12576 3120 12593 3184
rect 12657 3120 12674 3184
rect 12738 3120 12755 3184
rect 12819 3120 12836 3184
rect 12900 3120 12917 3184
rect 12981 3120 12998 3184
rect 13062 3120 13079 3184
rect 13143 3120 13160 3184
rect 13224 3120 13241 3184
rect 13305 3120 13322 3184
rect 13386 3120 13403 3184
rect 13467 3120 13484 3184
rect 13548 3120 13565 3184
rect 13629 3120 13646 3184
rect 13710 3120 13727 3184
rect 13791 3120 13808 3184
rect 13872 3120 13889 3184
rect 13953 3120 13970 3184
rect 14034 3120 14051 3184
rect 14115 3120 14132 3184
rect 14196 3120 14213 3184
rect 14277 3120 14294 3184
rect 14358 3120 14375 3184
rect 14439 3120 14456 3184
rect 14520 3120 14537 3184
rect 14601 3120 14618 3184
rect 14682 3120 14699 3184
rect 14763 3120 14780 3184
rect 14844 3120 14861 3184
rect 14925 3120 14931 3184
rect 10151 3096 14931 3120
rect 10151 3032 10157 3096
rect 10221 3032 10239 3096
rect 10303 3032 10321 3096
rect 10385 3032 10403 3096
rect 10467 3032 10485 3096
rect 10549 3032 10567 3096
rect 10631 3032 10649 3096
rect 10713 3032 10730 3096
rect 10794 3032 10811 3096
rect 10875 3032 10892 3096
rect 10956 3032 10973 3096
rect 11037 3032 11054 3096
rect 11118 3032 11135 3096
rect 11199 3032 11216 3096
rect 11280 3032 11297 3096
rect 11361 3032 11378 3096
rect 11442 3032 11459 3096
rect 11523 3032 11540 3096
rect 11604 3032 11621 3096
rect 11685 3032 11702 3096
rect 11766 3032 11783 3096
rect 11847 3032 11864 3096
rect 11928 3032 11945 3096
rect 12009 3032 12026 3096
rect 12090 3032 12107 3096
rect 12171 3032 12188 3096
rect 12252 3032 12269 3096
rect 12333 3032 12350 3096
rect 12414 3032 12431 3096
rect 12495 3032 12512 3096
rect 12576 3032 12593 3096
rect 12657 3032 12674 3096
rect 12738 3032 12755 3096
rect 12819 3032 12836 3096
rect 12900 3032 12917 3096
rect 12981 3032 12998 3096
rect 13062 3032 13079 3096
rect 13143 3032 13160 3096
rect 13224 3032 13241 3096
rect 13305 3032 13322 3096
rect 13386 3032 13403 3096
rect 13467 3032 13484 3096
rect 13548 3032 13565 3096
rect 13629 3032 13646 3096
rect 13710 3032 13727 3096
rect 13791 3032 13808 3096
rect 13872 3032 13889 3096
rect 13953 3032 13970 3096
rect 14034 3032 14051 3096
rect 14115 3032 14132 3096
rect 14196 3032 14213 3096
rect 14277 3032 14294 3096
rect 14358 3032 14375 3096
rect 14439 3032 14456 3096
rect 14520 3032 14537 3096
rect 14601 3032 14618 3096
rect 14682 3032 14699 3096
rect 14763 3032 14780 3096
rect 14844 3032 14861 3096
rect 14925 3032 14931 3096
rect 10151 3008 14931 3032
rect 10151 2944 10157 3008
rect 10221 2944 10239 3008
rect 10303 2944 10321 3008
rect 10385 2944 10403 3008
rect 10467 2944 10485 3008
rect 10549 2944 10567 3008
rect 10631 2944 10649 3008
rect 10713 2944 10730 3008
rect 10794 2944 10811 3008
rect 10875 2944 10892 3008
rect 10956 2944 10973 3008
rect 11037 2944 11054 3008
rect 11118 2944 11135 3008
rect 11199 2944 11216 3008
rect 11280 2944 11297 3008
rect 11361 2944 11378 3008
rect 11442 2944 11459 3008
rect 11523 2944 11540 3008
rect 11604 2944 11621 3008
rect 11685 2944 11702 3008
rect 11766 2944 11783 3008
rect 11847 2944 11864 3008
rect 11928 2944 11945 3008
rect 12009 2944 12026 3008
rect 12090 2944 12107 3008
rect 12171 2944 12188 3008
rect 12252 2944 12269 3008
rect 12333 2944 12350 3008
rect 12414 2944 12431 3008
rect 12495 2944 12512 3008
rect 12576 2944 12593 3008
rect 12657 2944 12674 3008
rect 12738 2944 12755 3008
rect 12819 2944 12836 3008
rect 12900 2944 12917 3008
rect 12981 2944 12998 3008
rect 13062 2944 13079 3008
rect 13143 2944 13160 3008
rect 13224 2944 13241 3008
rect 13305 2944 13322 3008
rect 13386 2944 13403 3008
rect 13467 2944 13484 3008
rect 13548 2944 13565 3008
rect 13629 2944 13646 3008
rect 13710 2944 13727 3008
rect 13791 2944 13808 3008
rect 13872 2944 13889 3008
rect 13953 2944 13970 3008
rect 14034 2944 14051 3008
rect 14115 2944 14132 3008
rect 14196 2944 14213 3008
rect 14277 2944 14294 3008
rect 14358 2944 14375 3008
rect 14439 2944 14456 3008
rect 14520 2944 14537 3008
rect 14601 2944 14618 3008
rect 14682 2944 14699 3008
rect 14763 2944 14780 3008
rect 14844 2944 14861 3008
rect 14925 2944 14931 3008
rect 10151 2920 14931 2944
rect 10151 2856 10157 2920
rect 10221 2856 10239 2920
rect 10303 2856 10321 2920
rect 10385 2856 10403 2920
rect 10467 2856 10485 2920
rect 10549 2856 10567 2920
rect 10631 2856 10649 2920
rect 10713 2856 10730 2920
rect 10794 2856 10811 2920
rect 10875 2856 10892 2920
rect 10956 2856 10973 2920
rect 11037 2856 11054 2920
rect 11118 2856 11135 2920
rect 11199 2856 11216 2920
rect 11280 2856 11297 2920
rect 11361 2856 11378 2920
rect 11442 2856 11459 2920
rect 11523 2856 11540 2920
rect 11604 2856 11621 2920
rect 11685 2856 11702 2920
rect 11766 2856 11783 2920
rect 11847 2856 11864 2920
rect 11928 2856 11945 2920
rect 12009 2856 12026 2920
rect 12090 2856 12107 2920
rect 12171 2856 12188 2920
rect 12252 2856 12269 2920
rect 12333 2856 12350 2920
rect 12414 2856 12431 2920
rect 12495 2856 12512 2920
rect 12576 2856 12593 2920
rect 12657 2856 12674 2920
rect 12738 2856 12755 2920
rect 12819 2856 12836 2920
rect 12900 2856 12917 2920
rect 12981 2856 12998 2920
rect 13062 2856 13079 2920
rect 13143 2856 13160 2920
rect 13224 2856 13241 2920
rect 13305 2856 13322 2920
rect 13386 2856 13403 2920
rect 13467 2856 13484 2920
rect 13548 2856 13565 2920
rect 13629 2856 13646 2920
rect 13710 2856 13727 2920
rect 13791 2856 13808 2920
rect 13872 2856 13889 2920
rect 13953 2856 13970 2920
rect 14034 2856 14051 2920
rect 14115 2856 14132 2920
rect 14196 2856 14213 2920
rect 14277 2856 14294 2920
rect 14358 2856 14375 2920
rect 14439 2856 14456 2920
rect 14520 2856 14537 2920
rect 14601 2856 14618 2920
rect 14682 2856 14699 2920
rect 14763 2856 14780 2920
rect 14844 2856 14861 2920
rect 14925 2856 14931 2920
rect 10151 2832 14931 2856
rect 10151 2768 10157 2832
rect 10221 2768 10239 2832
rect 10303 2768 10321 2832
rect 10385 2768 10403 2832
rect 10467 2768 10485 2832
rect 10549 2768 10567 2832
rect 10631 2768 10649 2832
rect 10713 2768 10730 2832
rect 10794 2768 10811 2832
rect 10875 2768 10892 2832
rect 10956 2768 10973 2832
rect 11037 2768 11054 2832
rect 11118 2768 11135 2832
rect 11199 2768 11216 2832
rect 11280 2768 11297 2832
rect 11361 2768 11378 2832
rect 11442 2768 11459 2832
rect 11523 2768 11540 2832
rect 11604 2768 11621 2832
rect 11685 2768 11702 2832
rect 11766 2768 11783 2832
rect 11847 2768 11864 2832
rect 11928 2768 11945 2832
rect 12009 2768 12026 2832
rect 12090 2768 12107 2832
rect 12171 2768 12188 2832
rect 12252 2768 12269 2832
rect 12333 2768 12350 2832
rect 12414 2768 12431 2832
rect 12495 2768 12512 2832
rect 12576 2768 12593 2832
rect 12657 2768 12674 2832
rect 12738 2768 12755 2832
rect 12819 2768 12836 2832
rect 12900 2768 12917 2832
rect 12981 2768 12998 2832
rect 13062 2768 13079 2832
rect 13143 2768 13160 2832
rect 13224 2768 13241 2832
rect 13305 2768 13322 2832
rect 13386 2768 13403 2832
rect 13467 2768 13484 2832
rect 13548 2768 13565 2832
rect 13629 2768 13646 2832
rect 13710 2768 13727 2832
rect 13791 2768 13808 2832
rect 13872 2768 13889 2832
rect 13953 2768 13970 2832
rect 14034 2768 14051 2832
rect 14115 2768 14132 2832
rect 14196 2768 14213 2832
rect 14277 2768 14294 2832
rect 14358 2768 14375 2832
rect 14439 2768 14456 2832
rect 14520 2768 14537 2832
rect 14601 2768 14618 2832
rect 14682 2768 14699 2832
rect 14763 2768 14780 2832
rect 14844 2768 14861 2832
rect 14925 2768 14931 2832
rect 10151 2744 14931 2768
rect 10151 2680 10157 2744
rect 10221 2680 10239 2744
rect 10303 2680 10321 2744
rect 10385 2680 10403 2744
rect 10467 2680 10485 2744
rect 10549 2680 10567 2744
rect 10631 2680 10649 2744
rect 10713 2680 10730 2744
rect 10794 2680 10811 2744
rect 10875 2680 10892 2744
rect 10956 2680 10973 2744
rect 11037 2680 11054 2744
rect 11118 2680 11135 2744
rect 11199 2680 11216 2744
rect 11280 2680 11297 2744
rect 11361 2680 11378 2744
rect 11442 2680 11459 2744
rect 11523 2680 11540 2744
rect 11604 2680 11621 2744
rect 11685 2680 11702 2744
rect 11766 2680 11783 2744
rect 11847 2680 11864 2744
rect 11928 2680 11945 2744
rect 12009 2680 12026 2744
rect 12090 2680 12107 2744
rect 12171 2680 12188 2744
rect 12252 2680 12269 2744
rect 12333 2680 12350 2744
rect 12414 2680 12431 2744
rect 12495 2680 12512 2744
rect 12576 2680 12593 2744
rect 12657 2680 12674 2744
rect 12738 2680 12755 2744
rect 12819 2680 12836 2744
rect 12900 2680 12917 2744
rect 12981 2680 12998 2744
rect 13062 2680 13079 2744
rect 13143 2680 13160 2744
rect 13224 2680 13241 2744
rect 13305 2680 13322 2744
rect 13386 2680 13403 2744
rect 13467 2680 13484 2744
rect 13548 2680 13565 2744
rect 13629 2680 13646 2744
rect 13710 2680 13727 2744
rect 13791 2680 13808 2744
rect 13872 2680 13889 2744
rect 13953 2680 13970 2744
rect 14034 2680 14051 2744
rect 14115 2680 14132 2744
rect 14196 2680 14213 2744
rect 14277 2680 14294 2744
rect 14358 2680 14375 2744
rect 14439 2680 14456 2744
rect 14520 2680 14537 2744
rect 14601 2680 14618 2744
rect 14682 2680 14699 2744
rect 14763 2680 14780 2744
rect 14844 2680 14861 2744
rect 14925 2680 14931 2744
rect 10151 2656 14931 2680
rect 10151 2592 10157 2656
rect 10221 2592 10239 2656
rect 10303 2592 10321 2656
rect 10385 2592 10403 2656
rect 10467 2592 10485 2656
rect 10549 2592 10567 2656
rect 10631 2592 10649 2656
rect 10713 2592 10730 2656
rect 10794 2592 10811 2656
rect 10875 2592 10892 2656
rect 10956 2592 10973 2656
rect 11037 2592 11054 2656
rect 11118 2592 11135 2656
rect 11199 2592 11216 2656
rect 11280 2592 11297 2656
rect 11361 2592 11378 2656
rect 11442 2592 11459 2656
rect 11523 2592 11540 2656
rect 11604 2592 11621 2656
rect 11685 2592 11702 2656
rect 11766 2592 11783 2656
rect 11847 2592 11864 2656
rect 11928 2592 11945 2656
rect 12009 2592 12026 2656
rect 12090 2592 12107 2656
rect 12171 2592 12188 2656
rect 12252 2592 12269 2656
rect 12333 2592 12350 2656
rect 12414 2592 12431 2656
rect 12495 2592 12512 2656
rect 12576 2592 12593 2656
rect 12657 2592 12674 2656
rect 12738 2592 12755 2656
rect 12819 2592 12836 2656
rect 12900 2592 12917 2656
rect 12981 2592 12998 2656
rect 13062 2592 13079 2656
rect 13143 2592 13160 2656
rect 13224 2592 13241 2656
rect 13305 2592 13322 2656
rect 13386 2592 13403 2656
rect 13467 2592 13484 2656
rect 13548 2592 13565 2656
rect 13629 2592 13646 2656
rect 13710 2592 13727 2656
rect 13791 2592 13808 2656
rect 13872 2592 13889 2656
rect 13953 2592 13970 2656
rect 14034 2592 14051 2656
rect 14115 2592 14132 2656
rect 14196 2592 14213 2656
rect 14277 2592 14294 2656
rect 14358 2592 14375 2656
rect 14439 2592 14456 2656
rect 14520 2592 14537 2656
rect 14601 2592 14618 2656
rect 14682 2592 14699 2656
rect 14763 2592 14780 2656
rect 14844 2592 14861 2656
rect 14925 2592 14931 2656
rect 10151 2588 14931 2592
<< via3 >>
rect 126 3208 190 3272
rect 208 3208 272 3272
rect 290 3208 354 3272
rect 372 3208 436 3272
rect 454 3208 518 3272
rect 536 3208 600 3272
rect 618 3208 682 3272
rect 699 3208 763 3272
rect 780 3208 844 3272
rect 861 3208 925 3272
rect 942 3208 1006 3272
rect 1023 3208 1087 3272
rect 1104 3208 1168 3272
rect 1185 3208 1249 3272
rect 1266 3208 1330 3272
rect 1347 3208 1411 3272
rect 1428 3208 1492 3272
rect 1509 3208 1573 3272
rect 1590 3208 1654 3272
rect 1671 3208 1735 3272
rect 1752 3208 1816 3272
rect 1833 3208 1897 3272
rect 1914 3208 1978 3272
rect 1995 3208 2059 3272
rect 2076 3208 2140 3272
rect 2157 3208 2221 3272
rect 2238 3208 2302 3272
rect 2319 3208 2383 3272
rect 2400 3208 2464 3272
rect 2481 3208 2545 3272
rect 2562 3208 2626 3272
rect 2643 3208 2707 3272
rect 2724 3208 2788 3272
rect 2805 3208 2869 3272
rect 2886 3208 2950 3272
rect 2967 3208 3031 3272
rect 3048 3208 3112 3272
rect 3129 3208 3193 3272
rect 3210 3208 3274 3272
rect 3291 3208 3355 3272
rect 3372 3208 3436 3272
rect 3453 3208 3517 3272
rect 3534 3208 3598 3272
rect 3615 3208 3679 3272
rect 3696 3208 3760 3272
rect 3777 3208 3841 3272
rect 3858 3208 3922 3272
rect 3939 3208 4003 3272
rect 4020 3208 4084 3272
rect 4101 3208 4165 3272
rect 4182 3208 4246 3272
rect 4263 3208 4327 3272
rect 4344 3208 4408 3272
rect 4425 3208 4489 3272
rect 4506 3208 4570 3272
rect 4587 3208 4651 3272
rect 4668 3208 4732 3272
rect 4749 3208 4813 3272
rect 4830 3208 4894 3272
rect 126 3120 190 3184
rect 208 3120 272 3184
rect 290 3120 354 3184
rect 372 3120 436 3184
rect 454 3120 518 3184
rect 536 3120 600 3184
rect 618 3120 682 3184
rect 699 3120 763 3184
rect 780 3120 844 3184
rect 861 3120 925 3184
rect 942 3120 1006 3184
rect 1023 3120 1087 3184
rect 1104 3120 1168 3184
rect 1185 3120 1249 3184
rect 1266 3120 1330 3184
rect 1347 3120 1411 3184
rect 1428 3120 1492 3184
rect 1509 3120 1573 3184
rect 1590 3120 1654 3184
rect 1671 3120 1735 3184
rect 1752 3120 1816 3184
rect 1833 3120 1897 3184
rect 1914 3120 1978 3184
rect 1995 3120 2059 3184
rect 2076 3120 2140 3184
rect 2157 3120 2221 3184
rect 2238 3120 2302 3184
rect 2319 3120 2383 3184
rect 2400 3120 2464 3184
rect 2481 3120 2545 3184
rect 2562 3120 2626 3184
rect 2643 3120 2707 3184
rect 2724 3120 2788 3184
rect 2805 3120 2869 3184
rect 2886 3120 2950 3184
rect 2967 3120 3031 3184
rect 3048 3120 3112 3184
rect 3129 3120 3193 3184
rect 3210 3120 3274 3184
rect 3291 3120 3355 3184
rect 3372 3120 3436 3184
rect 3453 3120 3517 3184
rect 3534 3120 3598 3184
rect 3615 3120 3679 3184
rect 3696 3120 3760 3184
rect 3777 3120 3841 3184
rect 3858 3120 3922 3184
rect 3939 3120 4003 3184
rect 4020 3120 4084 3184
rect 4101 3120 4165 3184
rect 4182 3120 4246 3184
rect 4263 3120 4327 3184
rect 4344 3120 4408 3184
rect 4425 3120 4489 3184
rect 4506 3120 4570 3184
rect 4587 3120 4651 3184
rect 4668 3120 4732 3184
rect 4749 3120 4813 3184
rect 4830 3120 4894 3184
rect 126 3032 190 3096
rect 208 3032 272 3096
rect 290 3032 354 3096
rect 372 3032 436 3096
rect 454 3032 518 3096
rect 536 3032 600 3096
rect 618 3032 682 3096
rect 699 3032 763 3096
rect 780 3032 844 3096
rect 861 3032 925 3096
rect 942 3032 1006 3096
rect 1023 3032 1087 3096
rect 1104 3032 1168 3096
rect 1185 3032 1249 3096
rect 1266 3032 1330 3096
rect 1347 3032 1411 3096
rect 1428 3032 1492 3096
rect 1509 3032 1573 3096
rect 1590 3032 1654 3096
rect 1671 3032 1735 3096
rect 1752 3032 1816 3096
rect 1833 3032 1897 3096
rect 1914 3032 1978 3096
rect 1995 3032 2059 3096
rect 2076 3032 2140 3096
rect 2157 3032 2221 3096
rect 2238 3032 2302 3096
rect 2319 3032 2383 3096
rect 2400 3032 2464 3096
rect 2481 3032 2545 3096
rect 2562 3032 2626 3096
rect 2643 3032 2707 3096
rect 2724 3032 2788 3096
rect 2805 3032 2869 3096
rect 2886 3032 2950 3096
rect 2967 3032 3031 3096
rect 3048 3032 3112 3096
rect 3129 3032 3193 3096
rect 3210 3032 3274 3096
rect 3291 3032 3355 3096
rect 3372 3032 3436 3096
rect 3453 3032 3517 3096
rect 3534 3032 3598 3096
rect 3615 3032 3679 3096
rect 3696 3032 3760 3096
rect 3777 3032 3841 3096
rect 3858 3032 3922 3096
rect 3939 3032 4003 3096
rect 4020 3032 4084 3096
rect 4101 3032 4165 3096
rect 4182 3032 4246 3096
rect 4263 3032 4327 3096
rect 4344 3032 4408 3096
rect 4425 3032 4489 3096
rect 4506 3032 4570 3096
rect 4587 3032 4651 3096
rect 4668 3032 4732 3096
rect 4749 3032 4813 3096
rect 4830 3032 4894 3096
rect 126 2944 190 3008
rect 208 2944 272 3008
rect 290 2944 354 3008
rect 372 2944 436 3008
rect 454 2944 518 3008
rect 536 2944 600 3008
rect 618 2944 682 3008
rect 699 2944 763 3008
rect 780 2944 844 3008
rect 861 2944 925 3008
rect 942 2944 1006 3008
rect 1023 2944 1087 3008
rect 1104 2944 1168 3008
rect 1185 2944 1249 3008
rect 1266 2944 1330 3008
rect 1347 2944 1411 3008
rect 1428 2944 1492 3008
rect 1509 2944 1573 3008
rect 1590 2944 1654 3008
rect 1671 2944 1735 3008
rect 1752 2944 1816 3008
rect 1833 2944 1897 3008
rect 1914 2944 1978 3008
rect 1995 2944 2059 3008
rect 2076 2944 2140 3008
rect 2157 2944 2221 3008
rect 2238 2944 2302 3008
rect 2319 2944 2383 3008
rect 2400 2944 2464 3008
rect 2481 2944 2545 3008
rect 2562 2944 2626 3008
rect 2643 2944 2707 3008
rect 2724 2944 2788 3008
rect 2805 2944 2869 3008
rect 2886 2944 2950 3008
rect 2967 2944 3031 3008
rect 3048 2944 3112 3008
rect 3129 2944 3193 3008
rect 3210 2944 3274 3008
rect 3291 2944 3355 3008
rect 3372 2944 3436 3008
rect 3453 2944 3517 3008
rect 3534 2944 3598 3008
rect 3615 2944 3679 3008
rect 3696 2944 3760 3008
rect 3777 2944 3841 3008
rect 3858 2944 3922 3008
rect 3939 2944 4003 3008
rect 4020 2944 4084 3008
rect 4101 2944 4165 3008
rect 4182 2944 4246 3008
rect 4263 2944 4327 3008
rect 4344 2944 4408 3008
rect 4425 2944 4489 3008
rect 4506 2944 4570 3008
rect 4587 2944 4651 3008
rect 4668 2944 4732 3008
rect 4749 2944 4813 3008
rect 4830 2944 4894 3008
rect 126 2856 190 2920
rect 208 2856 272 2920
rect 290 2856 354 2920
rect 372 2856 436 2920
rect 454 2856 518 2920
rect 536 2856 600 2920
rect 618 2856 682 2920
rect 699 2856 763 2920
rect 780 2856 844 2920
rect 861 2856 925 2920
rect 942 2856 1006 2920
rect 1023 2856 1087 2920
rect 1104 2856 1168 2920
rect 1185 2856 1249 2920
rect 1266 2856 1330 2920
rect 1347 2856 1411 2920
rect 1428 2856 1492 2920
rect 1509 2856 1573 2920
rect 1590 2856 1654 2920
rect 1671 2856 1735 2920
rect 1752 2856 1816 2920
rect 1833 2856 1897 2920
rect 1914 2856 1978 2920
rect 1995 2856 2059 2920
rect 2076 2856 2140 2920
rect 2157 2856 2221 2920
rect 2238 2856 2302 2920
rect 2319 2856 2383 2920
rect 2400 2856 2464 2920
rect 2481 2856 2545 2920
rect 2562 2856 2626 2920
rect 2643 2856 2707 2920
rect 2724 2856 2788 2920
rect 2805 2856 2869 2920
rect 2886 2856 2950 2920
rect 2967 2856 3031 2920
rect 3048 2856 3112 2920
rect 3129 2856 3193 2920
rect 3210 2856 3274 2920
rect 3291 2856 3355 2920
rect 3372 2856 3436 2920
rect 3453 2856 3517 2920
rect 3534 2856 3598 2920
rect 3615 2856 3679 2920
rect 3696 2856 3760 2920
rect 3777 2856 3841 2920
rect 3858 2856 3922 2920
rect 3939 2856 4003 2920
rect 4020 2856 4084 2920
rect 4101 2856 4165 2920
rect 4182 2856 4246 2920
rect 4263 2856 4327 2920
rect 4344 2856 4408 2920
rect 4425 2856 4489 2920
rect 4506 2856 4570 2920
rect 4587 2856 4651 2920
rect 4668 2856 4732 2920
rect 4749 2856 4813 2920
rect 4830 2856 4894 2920
rect 126 2768 190 2832
rect 208 2768 272 2832
rect 290 2768 354 2832
rect 372 2768 436 2832
rect 454 2768 518 2832
rect 536 2768 600 2832
rect 618 2768 682 2832
rect 699 2768 763 2832
rect 780 2768 844 2832
rect 861 2768 925 2832
rect 942 2768 1006 2832
rect 1023 2768 1087 2832
rect 1104 2768 1168 2832
rect 1185 2768 1249 2832
rect 1266 2768 1330 2832
rect 1347 2768 1411 2832
rect 1428 2768 1492 2832
rect 1509 2768 1573 2832
rect 1590 2768 1654 2832
rect 1671 2768 1735 2832
rect 1752 2768 1816 2832
rect 1833 2768 1897 2832
rect 1914 2768 1978 2832
rect 1995 2768 2059 2832
rect 2076 2768 2140 2832
rect 2157 2768 2221 2832
rect 2238 2768 2302 2832
rect 2319 2768 2383 2832
rect 2400 2768 2464 2832
rect 2481 2768 2545 2832
rect 2562 2768 2626 2832
rect 2643 2768 2707 2832
rect 2724 2768 2788 2832
rect 2805 2768 2869 2832
rect 2886 2768 2950 2832
rect 2967 2768 3031 2832
rect 3048 2768 3112 2832
rect 3129 2768 3193 2832
rect 3210 2768 3274 2832
rect 3291 2768 3355 2832
rect 3372 2768 3436 2832
rect 3453 2768 3517 2832
rect 3534 2768 3598 2832
rect 3615 2768 3679 2832
rect 3696 2768 3760 2832
rect 3777 2768 3841 2832
rect 3858 2768 3922 2832
rect 3939 2768 4003 2832
rect 4020 2768 4084 2832
rect 4101 2768 4165 2832
rect 4182 2768 4246 2832
rect 4263 2768 4327 2832
rect 4344 2768 4408 2832
rect 4425 2768 4489 2832
rect 4506 2768 4570 2832
rect 4587 2768 4651 2832
rect 4668 2768 4732 2832
rect 4749 2768 4813 2832
rect 4830 2768 4894 2832
rect 126 2680 190 2744
rect 208 2680 272 2744
rect 290 2680 354 2744
rect 372 2680 436 2744
rect 454 2680 518 2744
rect 536 2680 600 2744
rect 618 2680 682 2744
rect 699 2680 763 2744
rect 780 2680 844 2744
rect 861 2680 925 2744
rect 942 2680 1006 2744
rect 1023 2680 1087 2744
rect 1104 2680 1168 2744
rect 1185 2680 1249 2744
rect 1266 2680 1330 2744
rect 1347 2680 1411 2744
rect 1428 2680 1492 2744
rect 1509 2680 1573 2744
rect 1590 2680 1654 2744
rect 1671 2680 1735 2744
rect 1752 2680 1816 2744
rect 1833 2680 1897 2744
rect 1914 2680 1978 2744
rect 1995 2680 2059 2744
rect 2076 2680 2140 2744
rect 2157 2680 2221 2744
rect 2238 2680 2302 2744
rect 2319 2680 2383 2744
rect 2400 2680 2464 2744
rect 2481 2680 2545 2744
rect 2562 2680 2626 2744
rect 2643 2680 2707 2744
rect 2724 2680 2788 2744
rect 2805 2680 2869 2744
rect 2886 2680 2950 2744
rect 2967 2680 3031 2744
rect 3048 2680 3112 2744
rect 3129 2680 3193 2744
rect 3210 2680 3274 2744
rect 3291 2680 3355 2744
rect 3372 2680 3436 2744
rect 3453 2680 3517 2744
rect 3534 2680 3598 2744
rect 3615 2680 3679 2744
rect 3696 2680 3760 2744
rect 3777 2680 3841 2744
rect 3858 2680 3922 2744
rect 3939 2680 4003 2744
rect 4020 2680 4084 2744
rect 4101 2680 4165 2744
rect 4182 2680 4246 2744
rect 4263 2680 4327 2744
rect 4344 2680 4408 2744
rect 4425 2680 4489 2744
rect 4506 2680 4570 2744
rect 4587 2680 4651 2744
rect 4668 2680 4732 2744
rect 4749 2680 4813 2744
rect 4830 2680 4894 2744
rect 126 2592 190 2656
rect 208 2592 272 2656
rect 290 2592 354 2656
rect 372 2592 436 2656
rect 454 2592 518 2656
rect 536 2592 600 2656
rect 618 2592 682 2656
rect 699 2592 763 2656
rect 780 2592 844 2656
rect 861 2592 925 2656
rect 942 2592 1006 2656
rect 1023 2592 1087 2656
rect 1104 2592 1168 2656
rect 1185 2592 1249 2656
rect 1266 2592 1330 2656
rect 1347 2592 1411 2656
rect 1428 2592 1492 2656
rect 1509 2592 1573 2656
rect 1590 2592 1654 2656
rect 1671 2592 1735 2656
rect 1752 2592 1816 2656
rect 1833 2592 1897 2656
rect 1914 2592 1978 2656
rect 1995 2592 2059 2656
rect 2076 2592 2140 2656
rect 2157 2592 2221 2656
rect 2238 2592 2302 2656
rect 2319 2592 2383 2656
rect 2400 2592 2464 2656
rect 2481 2592 2545 2656
rect 2562 2592 2626 2656
rect 2643 2592 2707 2656
rect 2724 2592 2788 2656
rect 2805 2592 2869 2656
rect 2886 2592 2950 2656
rect 2967 2592 3031 2656
rect 3048 2592 3112 2656
rect 3129 2592 3193 2656
rect 3210 2592 3274 2656
rect 3291 2592 3355 2656
rect 3372 2592 3436 2656
rect 3453 2592 3517 2656
rect 3534 2592 3598 2656
rect 3615 2592 3679 2656
rect 3696 2592 3760 2656
rect 3777 2592 3841 2656
rect 3858 2592 3922 2656
rect 3939 2592 4003 2656
rect 4020 2592 4084 2656
rect 4101 2592 4165 2656
rect 4182 2592 4246 2656
rect 4263 2592 4327 2656
rect 4344 2592 4408 2656
rect 4425 2592 4489 2656
rect 4506 2592 4570 2656
rect 4587 2592 4651 2656
rect 4668 2592 4732 2656
rect 4749 2592 4813 2656
rect 4830 2592 4894 2656
rect 10157 3208 10221 3272
rect 10239 3208 10303 3272
rect 10321 3208 10385 3272
rect 10403 3208 10467 3272
rect 10485 3208 10549 3272
rect 10567 3208 10631 3272
rect 10649 3208 10713 3272
rect 10730 3208 10794 3272
rect 10811 3208 10875 3272
rect 10892 3208 10956 3272
rect 10973 3208 11037 3272
rect 11054 3208 11118 3272
rect 11135 3208 11199 3272
rect 11216 3208 11280 3272
rect 11297 3208 11361 3272
rect 11378 3208 11442 3272
rect 11459 3208 11523 3272
rect 11540 3208 11604 3272
rect 11621 3208 11685 3272
rect 11702 3208 11766 3272
rect 11783 3208 11847 3272
rect 11864 3208 11928 3272
rect 11945 3208 12009 3272
rect 12026 3208 12090 3272
rect 12107 3208 12171 3272
rect 12188 3208 12252 3272
rect 12269 3208 12333 3272
rect 12350 3208 12414 3272
rect 12431 3208 12495 3272
rect 12512 3208 12576 3272
rect 12593 3208 12657 3272
rect 12674 3208 12738 3272
rect 12755 3208 12819 3272
rect 12836 3208 12900 3272
rect 12917 3208 12981 3272
rect 12998 3208 13062 3272
rect 13079 3208 13143 3272
rect 13160 3208 13224 3272
rect 13241 3208 13305 3272
rect 13322 3208 13386 3272
rect 13403 3208 13467 3272
rect 13484 3208 13548 3272
rect 13565 3208 13629 3272
rect 13646 3208 13710 3272
rect 13727 3208 13791 3272
rect 13808 3208 13872 3272
rect 13889 3208 13953 3272
rect 13970 3208 14034 3272
rect 14051 3208 14115 3272
rect 14132 3208 14196 3272
rect 14213 3208 14277 3272
rect 14294 3208 14358 3272
rect 14375 3208 14439 3272
rect 14456 3208 14520 3272
rect 14537 3208 14601 3272
rect 14618 3208 14682 3272
rect 14699 3208 14763 3272
rect 14780 3208 14844 3272
rect 14861 3208 14925 3272
rect 10157 3120 10221 3184
rect 10239 3120 10303 3184
rect 10321 3120 10385 3184
rect 10403 3120 10467 3184
rect 10485 3120 10549 3184
rect 10567 3120 10631 3184
rect 10649 3120 10713 3184
rect 10730 3120 10794 3184
rect 10811 3120 10875 3184
rect 10892 3120 10956 3184
rect 10973 3120 11037 3184
rect 11054 3120 11118 3184
rect 11135 3120 11199 3184
rect 11216 3120 11280 3184
rect 11297 3120 11361 3184
rect 11378 3120 11442 3184
rect 11459 3120 11523 3184
rect 11540 3120 11604 3184
rect 11621 3120 11685 3184
rect 11702 3120 11766 3184
rect 11783 3120 11847 3184
rect 11864 3120 11928 3184
rect 11945 3120 12009 3184
rect 12026 3120 12090 3184
rect 12107 3120 12171 3184
rect 12188 3120 12252 3184
rect 12269 3120 12333 3184
rect 12350 3120 12414 3184
rect 12431 3120 12495 3184
rect 12512 3120 12576 3184
rect 12593 3120 12657 3184
rect 12674 3120 12738 3184
rect 12755 3120 12819 3184
rect 12836 3120 12900 3184
rect 12917 3120 12981 3184
rect 12998 3120 13062 3184
rect 13079 3120 13143 3184
rect 13160 3120 13224 3184
rect 13241 3120 13305 3184
rect 13322 3120 13386 3184
rect 13403 3120 13467 3184
rect 13484 3120 13548 3184
rect 13565 3120 13629 3184
rect 13646 3120 13710 3184
rect 13727 3120 13791 3184
rect 13808 3120 13872 3184
rect 13889 3120 13953 3184
rect 13970 3120 14034 3184
rect 14051 3120 14115 3184
rect 14132 3120 14196 3184
rect 14213 3120 14277 3184
rect 14294 3120 14358 3184
rect 14375 3120 14439 3184
rect 14456 3120 14520 3184
rect 14537 3120 14601 3184
rect 14618 3120 14682 3184
rect 14699 3120 14763 3184
rect 14780 3120 14844 3184
rect 14861 3120 14925 3184
rect 10157 3032 10221 3096
rect 10239 3032 10303 3096
rect 10321 3032 10385 3096
rect 10403 3032 10467 3096
rect 10485 3032 10549 3096
rect 10567 3032 10631 3096
rect 10649 3032 10713 3096
rect 10730 3032 10794 3096
rect 10811 3032 10875 3096
rect 10892 3032 10956 3096
rect 10973 3032 11037 3096
rect 11054 3032 11118 3096
rect 11135 3032 11199 3096
rect 11216 3032 11280 3096
rect 11297 3032 11361 3096
rect 11378 3032 11442 3096
rect 11459 3032 11523 3096
rect 11540 3032 11604 3096
rect 11621 3032 11685 3096
rect 11702 3032 11766 3096
rect 11783 3032 11847 3096
rect 11864 3032 11928 3096
rect 11945 3032 12009 3096
rect 12026 3032 12090 3096
rect 12107 3032 12171 3096
rect 12188 3032 12252 3096
rect 12269 3032 12333 3096
rect 12350 3032 12414 3096
rect 12431 3032 12495 3096
rect 12512 3032 12576 3096
rect 12593 3032 12657 3096
rect 12674 3032 12738 3096
rect 12755 3032 12819 3096
rect 12836 3032 12900 3096
rect 12917 3032 12981 3096
rect 12998 3032 13062 3096
rect 13079 3032 13143 3096
rect 13160 3032 13224 3096
rect 13241 3032 13305 3096
rect 13322 3032 13386 3096
rect 13403 3032 13467 3096
rect 13484 3032 13548 3096
rect 13565 3032 13629 3096
rect 13646 3032 13710 3096
rect 13727 3032 13791 3096
rect 13808 3032 13872 3096
rect 13889 3032 13953 3096
rect 13970 3032 14034 3096
rect 14051 3032 14115 3096
rect 14132 3032 14196 3096
rect 14213 3032 14277 3096
rect 14294 3032 14358 3096
rect 14375 3032 14439 3096
rect 14456 3032 14520 3096
rect 14537 3032 14601 3096
rect 14618 3032 14682 3096
rect 14699 3032 14763 3096
rect 14780 3032 14844 3096
rect 14861 3032 14925 3096
rect 10157 2944 10221 3008
rect 10239 2944 10303 3008
rect 10321 2944 10385 3008
rect 10403 2944 10467 3008
rect 10485 2944 10549 3008
rect 10567 2944 10631 3008
rect 10649 2944 10713 3008
rect 10730 2944 10794 3008
rect 10811 2944 10875 3008
rect 10892 2944 10956 3008
rect 10973 2944 11037 3008
rect 11054 2944 11118 3008
rect 11135 2944 11199 3008
rect 11216 2944 11280 3008
rect 11297 2944 11361 3008
rect 11378 2944 11442 3008
rect 11459 2944 11523 3008
rect 11540 2944 11604 3008
rect 11621 2944 11685 3008
rect 11702 2944 11766 3008
rect 11783 2944 11847 3008
rect 11864 2944 11928 3008
rect 11945 2944 12009 3008
rect 12026 2944 12090 3008
rect 12107 2944 12171 3008
rect 12188 2944 12252 3008
rect 12269 2944 12333 3008
rect 12350 2944 12414 3008
rect 12431 2944 12495 3008
rect 12512 2944 12576 3008
rect 12593 2944 12657 3008
rect 12674 2944 12738 3008
rect 12755 2944 12819 3008
rect 12836 2944 12900 3008
rect 12917 2944 12981 3008
rect 12998 2944 13062 3008
rect 13079 2944 13143 3008
rect 13160 2944 13224 3008
rect 13241 2944 13305 3008
rect 13322 2944 13386 3008
rect 13403 2944 13467 3008
rect 13484 2944 13548 3008
rect 13565 2944 13629 3008
rect 13646 2944 13710 3008
rect 13727 2944 13791 3008
rect 13808 2944 13872 3008
rect 13889 2944 13953 3008
rect 13970 2944 14034 3008
rect 14051 2944 14115 3008
rect 14132 2944 14196 3008
rect 14213 2944 14277 3008
rect 14294 2944 14358 3008
rect 14375 2944 14439 3008
rect 14456 2944 14520 3008
rect 14537 2944 14601 3008
rect 14618 2944 14682 3008
rect 14699 2944 14763 3008
rect 14780 2944 14844 3008
rect 14861 2944 14925 3008
rect 10157 2856 10221 2920
rect 10239 2856 10303 2920
rect 10321 2856 10385 2920
rect 10403 2856 10467 2920
rect 10485 2856 10549 2920
rect 10567 2856 10631 2920
rect 10649 2856 10713 2920
rect 10730 2856 10794 2920
rect 10811 2856 10875 2920
rect 10892 2856 10956 2920
rect 10973 2856 11037 2920
rect 11054 2856 11118 2920
rect 11135 2856 11199 2920
rect 11216 2856 11280 2920
rect 11297 2856 11361 2920
rect 11378 2856 11442 2920
rect 11459 2856 11523 2920
rect 11540 2856 11604 2920
rect 11621 2856 11685 2920
rect 11702 2856 11766 2920
rect 11783 2856 11847 2920
rect 11864 2856 11928 2920
rect 11945 2856 12009 2920
rect 12026 2856 12090 2920
rect 12107 2856 12171 2920
rect 12188 2856 12252 2920
rect 12269 2856 12333 2920
rect 12350 2856 12414 2920
rect 12431 2856 12495 2920
rect 12512 2856 12576 2920
rect 12593 2856 12657 2920
rect 12674 2856 12738 2920
rect 12755 2856 12819 2920
rect 12836 2856 12900 2920
rect 12917 2856 12981 2920
rect 12998 2856 13062 2920
rect 13079 2856 13143 2920
rect 13160 2856 13224 2920
rect 13241 2856 13305 2920
rect 13322 2856 13386 2920
rect 13403 2856 13467 2920
rect 13484 2856 13548 2920
rect 13565 2856 13629 2920
rect 13646 2856 13710 2920
rect 13727 2856 13791 2920
rect 13808 2856 13872 2920
rect 13889 2856 13953 2920
rect 13970 2856 14034 2920
rect 14051 2856 14115 2920
rect 14132 2856 14196 2920
rect 14213 2856 14277 2920
rect 14294 2856 14358 2920
rect 14375 2856 14439 2920
rect 14456 2856 14520 2920
rect 14537 2856 14601 2920
rect 14618 2856 14682 2920
rect 14699 2856 14763 2920
rect 14780 2856 14844 2920
rect 14861 2856 14925 2920
rect 10157 2768 10221 2832
rect 10239 2768 10303 2832
rect 10321 2768 10385 2832
rect 10403 2768 10467 2832
rect 10485 2768 10549 2832
rect 10567 2768 10631 2832
rect 10649 2768 10713 2832
rect 10730 2768 10794 2832
rect 10811 2768 10875 2832
rect 10892 2768 10956 2832
rect 10973 2768 11037 2832
rect 11054 2768 11118 2832
rect 11135 2768 11199 2832
rect 11216 2768 11280 2832
rect 11297 2768 11361 2832
rect 11378 2768 11442 2832
rect 11459 2768 11523 2832
rect 11540 2768 11604 2832
rect 11621 2768 11685 2832
rect 11702 2768 11766 2832
rect 11783 2768 11847 2832
rect 11864 2768 11928 2832
rect 11945 2768 12009 2832
rect 12026 2768 12090 2832
rect 12107 2768 12171 2832
rect 12188 2768 12252 2832
rect 12269 2768 12333 2832
rect 12350 2768 12414 2832
rect 12431 2768 12495 2832
rect 12512 2768 12576 2832
rect 12593 2768 12657 2832
rect 12674 2768 12738 2832
rect 12755 2768 12819 2832
rect 12836 2768 12900 2832
rect 12917 2768 12981 2832
rect 12998 2768 13062 2832
rect 13079 2768 13143 2832
rect 13160 2768 13224 2832
rect 13241 2768 13305 2832
rect 13322 2768 13386 2832
rect 13403 2768 13467 2832
rect 13484 2768 13548 2832
rect 13565 2768 13629 2832
rect 13646 2768 13710 2832
rect 13727 2768 13791 2832
rect 13808 2768 13872 2832
rect 13889 2768 13953 2832
rect 13970 2768 14034 2832
rect 14051 2768 14115 2832
rect 14132 2768 14196 2832
rect 14213 2768 14277 2832
rect 14294 2768 14358 2832
rect 14375 2768 14439 2832
rect 14456 2768 14520 2832
rect 14537 2768 14601 2832
rect 14618 2768 14682 2832
rect 14699 2768 14763 2832
rect 14780 2768 14844 2832
rect 14861 2768 14925 2832
rect 10157 2680 10221 2744
rect 10239 2680 10303 2744
rect 10321 2680 10385 2744
rect 10403 2680 10467 2744
rect 10485 2680 10549 2744
rect 10567 2680 10631 2744
rect 10649 2680 10713 2744
rect 10730 2680 10794 2744
rect 10811 2680 10875 2744
rect 10892 2680 10956 2744
rect 10973 2680 11037 2744
rect 11054 2680 11118 2744
rect 11135 2680 11199 2744
rect 11216 2680 11280 2744
rect 11297 2680 11361 2744
rect 11378 2680 11442 2744
rect 11459 2680 11523 2744
rect 11540 2680 11604 2744
rect 11621 2680 11685 2744
rect 11702 2680 11766 2744
rect 11783 2680 11847 2744
rect 11864 2680 11928 2744
rect 11945 2680 12009 2744
rect 12026 2680 12090 2744
rect 12107 2680 12171 2744
rect 12188 2680 12252 2744
rect 12269 2680 12333 2744
rect 12350 2680 12414 2744
rect 12431 2680 12495 2744
rect 12512 2680 12576 2744
rect 12593 2680 12657 2744
rect 12674 2680 12738 2744
rect 12755 2680 12819 2744
rect 12836 2680 12900 2744
rect 12917 2680 12981 2744
rect 12998 2680 13062 2744
rect 13079 2680 13143 2744
rect 13160 2680 13224 2744
rect 13241 2680 13305 2744
rect 13322 2680 13386 2744
rect 13403 2680 13467 2744
rect 13484 2680 13548 2744
rect 13565 2680 13629 2744
rect 13646 2680 13710 2744
rect 13727 2680 13791 2744
rect 13808 2680 13872 2744
rect 13889 2680 13953 2744
rect 13970 2680 14034 2744
rect 14051 2680 14115 2744
rect 14132 2680 14196 2744
rect 14213 2680 14277 2744
rect 14294 2680 14358 2744
rect 14375 2680 14439 2744
rect 14456 2680 14520 2744
rect 14537 2680 14601 2744
rect 14618 2680 14682 2744
rect 14699 2680 14763 2744
rect 14780 2680 14844 2744
rect 14861 2680 14925 2744
rect 10157 2592 10221 2656
rect 10239 2592 10303 2656
rect 10321 2592 10385 2656
rect 10403 2592 10467 2656
rect 10485 2592 10549 2656
rect 10567 2592 10631 2656
rect 10649 2592 10713 2656
rect 10730 2592 10794 2656
rect 10811 2592 10875 2656
rect 10892 2592 10956 2656
rect 10973 2592 11037 2656
rect 11054 2592 11118 2656
rect 11135 2592 11199 2656
rect 11216 2592 11280 2656
rect 11297 2592 11361 2656
rect 11378 2592 11442 2656
rect 11459 2592 11523 2656
rect 11540 2592 11604 2656
rect 11621 2592 11685 2656
rect 11702 2592 11766 2656
rect 11783 2592 11847 2656
rect 11864 2592 11928 2656
rect 11945 2592 12009 2656
rect 12026 2592 12090 2656
rect 12107 2592 12171 2656
rect 12188 2592 12252 2656
rect 12269 2592 12333 2656
rect 12350 2592 12414 2656
rect 12431 2592 12495 2656
rect 12512 2592 12576 2656
rect 12593 2592 12657 2656
rect 12674 2592 12738 2656
rect 12755 2592 12819 2656
rect 12836 2592 12900 2656
rect 12917 2592 12981 2656
rect 12998 2592 13062 2656
rect 13079 2592 13143 2656
rect 13160 2592 13224 2656
rect 13241 2592 13305 2656
rect 13322 2592 13386 2656
rect 13403 2592 13467 2656
rect 13484 2592 13548 2656
rect 13565 2592 13629 2656
rect 13646 2592 13710 2656
rect 13727 2592 13791 2656
rect 13808 2592 13872 2656
rect 13889 2592 13953 2656
rect 13970 2592 14034 2656
rect 14051 2592 14115 2656
rect 14132 2592 14196 2656
rect 14213 2592 14277 2656
rect 14294 2592 14358 2656
rect 14375 2592 14439 2656
rect 14456 2592 14520 2656
rect 14537 2592 14601 2656
rect 14618 2592 14682 2656
rect 14699 2592 14763 2656
rect 14780 2592 14844 2656
rect 14861 2592 14925 2656
<< metal4 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18600
rect 14746 13607 15000 18600
rect 0 12417 254 13307
rect 14746 12417 15000 13307
rect 0 11247 254 12137
rect 14746 11247 15000 12137
rect 0 10881 254 10947
rect 14746 10881 15000 10947
rect 0 10225 254 10821
rect 14746 10225 15000 10821
rect 0 9929 254 10165
rect 14746 9929 15000 10165
rect 0 9273 254 9869
rect 14746 9273 15000 9869
rect 0 9147 254 9213
rect 14746 9147 15000 9213
rect 0 7917 254 8847
rect 14746 7917 15000 8847
rect 0 6947 254 7637
rect 14746 6947 15000 7637
rect 0 5977 254 6667
rect 14746 5977 15000 6667
rect 0 4767 254 5697
rect 14746 4767 15000 5697
rect 0 3557 254 4487
rect 14746 3557 15000 4487
rect 0 3272 4895 3277
rect 0 3208 126 3272
rect 190 3208 208 3272
rect 272 3208 290 3272
rect 354 3208 372 3272
rect 436 3208 454 3272
rect 518 3208 536 3272
rect 600 3208 618 3272
rect 682 3208 699 3272
rect 763 3208 780 3272
rect 844 3208 861 3272
rect 925 3208 942 3272
rect 1006 3208 1023 3272
rect 1087 3208 1104 3272
rect 1168 3208 1185 3272
rect 1249 3208 1266 3272
rect 1330 3208 1347 3272
rect 1411 3208 1428 3272
rect 1492 3208 1509 3272
rect 1573 3208 1590 3272
rect 1654 3208 1671 3272
rect 1735 3208 1752 3272
rect 1816 3208 1833 3272
rect 1897 3208 1914 3272
rect 1978 3208 1995 3272
rect 2059 3208 2076 3272
rect 2140 3208 2157 3272
rect 2221 3208 2238 3272
rect 2302 3208 2319 3272
rect 2383 3208 2400 3272
rect 2464 3208 2481 3272
rect 2545 3208 2562 3272
rect 2626 3208 2643 3272
rect 2707 3208 2724 3272
rect 2788 3208 2805 3272
rect 2869 3208 2886 3272
rect 2950 3208 2967 3272
rect 3031 3208 3048 3272
rect 3112 3208 3129 3272
rect 3193 3208 3210 3272
rect 3274 3208 3291 3272
rect 3355 3208 3372 3272
rect 3436 3208 3453 3272
rect 3517 3208 3534 3272
rect 3598 3208 3615 3272
rect 3679 3208 3696 3272
rect 3760 3208 3777 3272
rect 3841 3208 3858 3272
rect 3922 3208 3939 3272
rect 4003 3208 4020 3272
rect 4084 3208 4101 3272
rect 4165 3208 4182 3272
rect 4246 3208 4263 3272
rect 4327 3208 4344 3272
rect 4408 3208 4425 3272
rect 4489 3208 4506 3272
rect 4570 3208 4587 3272
rect 4651 3208 4668 3272
rect 4732 3208 4749 3272
rect 4813 3208 4830 3272
rect 4894 3208 4895 3272
rect 0 3184 4895 3208
rect 0 3120 126 3184
rect 190 3120 208 3184
rect 272 3120 290 3184
rect 354 3120 372 3184
rect 436 3120 454 3184
rect 518 3120 536 3184
rect 600 3120 618 3184
rect 682 3120 699 3184
rect 763 3120 780 3184
rect 844 3120 861 3184
rect 925 3120 942 3184
rect 1006 3120 1023 3184
rect 1087 3120 1104 3184
rect 1168 3120 1185 3184
rect 1249 3120 1266 3184
rect 1330 3120 1347 3184
rect 1411 3120 1428 3184
rect 1492 3120 1509 3184
rect 1573 3120 1590 3184
rect 1654 3120 1671 3184
rect 1735 3120 1752 3184
rect 1816 3120 1833 3184
rect 1897 3120 1914 3184
rect 1978 3120 1995 3184
rect 2059 3120 2076 3184
rect 2140 3120 2157 3184
rect 2221 3120 2238 3184
rect 2302 3120 2319 3184
rect 2383 3120 2400 3184
rect 2464 3120 2481 3184
rect 2545 3120 2562 3184
rect 2626 3120 2643 3184
rect 2707 3120 2724 3184
rect 2788 3120 2805 3184
rect 2869 3120 2886 3184
rect 2950 3120 2967 3184
rect 3031 3120 3048 3184
rect 3112 3120 3129 3184
rect 3193 3120 3210 3184
rect 3274 3120 3291 3184
rect 3355 3120 3372 3184
rect 3436 3120 3453 3184
rect 3517 3120 3534 3184
rect 3598 3120 3615 3184
rect 3679 3120 3696 3184
rect 3760 3120 3777 3184
rect 3841 3120 3858 3184
rect 3922 3120 3939 3184
rect 4003 3120 4020 3184
rect 4084 3120 4101 3184
rect 4165 3120 4182 3184
rect 4246 3120 4263 3184
rect 4327 3120 4344 3184
rect 4408 3120 4425 3184
rect 4489 3120 4506 3184
rect 4570 3120 4587 3184
rect 4651 3120 4668 3184
rect 4732 3120 4749 3184
rect 4813 3120 4830 3184
rect 4894 3120 4895 3184
rect 0 3096 4895 3120
rect 0 3032 126 3096
rect 190 3032 208 3096
rect 272 3032 290 3096
rect 354 3032 372 3096
rect 436 3032 454 3096
rect 518 3032 536 3096
rect 600 3032 618 3096
rect 682 3032 699 3096
rect 763 3032 780 3096
rect 844 3032 861 3096
rect 925 3032 942 3096
rect 1006 3032 1023 3096
rect 1087 3032 1104 3096
rect 1168 3032 1185 3096
rect 1249 3032 1266 3096
rect 1330 3032 1347 3096
rect 1411 3032 1428 3096
rect 1492 3032 1509 3096
rect 1573 3032 1590 3096
rect 1654 3032 1671 3096
rect 1735 3032 1752 3096
rect 1816 3032 1833 3096
rect 1897 3032 1914 3096
rect 1978 3032 1995 3096
rect 2059 3032 2076 3096
rect 2140 3032 2157 3096
rect 2221 3032 2238 3096
rect 2302 3032 2319 3096
rect 2383 3032 2400 3096
rect 2464 3032 2481 3096
rect 2545 3032 2562 3096
rect 2626 3032 2643 3096
rect 2707 3032 2724 3096
rect 2788 3032 2805 3096
rect 2869 3032 2886 3096
rect 2950 3032 2967 3096
rect 3031 3032 3048 3096
rect 3112 3032 3129 3096
rect 3193 3032 3210 3096
rect 3274 3032 3291 3096
rect 3355 3032 3372 3096
rect 3436 3032 3453 3096
rect 3517 3032 3534 3096
rect 3598 3032 3615 3096
rect 3679 3032 3696 3096
rect 3760 3032 3777 3096
rect 3841 3032 3858 3096
rect 3922 3032 3939 3096
rect 4003 3032 4020 3096
rect 4084 3032 4101 3096
rect 4165 3032 4182 3096
rect 4246 3032 4263 3096
rect 4327 3032 4344 3096
rect 4408 3032 4425 3096
rect 4489 3032 4506 3096
rect 4570 3032 4587 3096
rect 4651 3032 4668 3096
rect 4732 3032 4749 3096
rect 4813 3032 4830 3096
rect 4894 3032 4895 3096
rect 0 3008 4895 3032
rect 0 2944 126 3008
rect 190 2944 208 3008
rect 272 2944 290 3008
rect 354 2944 372 3008
rect 436 2944 454 3008
rect 518 2944 536 3008
rect 600 2944 618 3008
rect 682 2944 699 3008
rect 763 2944 780 3008
rect 844 2944 861 3008
rect 925 2944 942 3008
rect 1006 2944 1023 3008
rect 1087 2944 1104 3008
rect 1168 2944 1185 3008
rect 1249 2944 1266 3008
rect 1330 2944 1347 3008
rect 1411 2944 1428 3008
rect 1492 2944 1509 3008
rect 1573 2944 1590 3008
rect 1654 2944 1671 3008
rect 1735 2944 1752 3008
rect 1816 2944 1833 3008
rect 1897 2944 1914 3008
rect 1978 2944 1995 3008
rect 2059 2944 2076 3008
rect 2140 2944 2157 3008
rect 2221 2944 2238 3008
rect 2302 2944 2319 3008
rect 2383 2944 2400 3008
rect 2464 2944 2481 3008
rect 2545 2944 2562 3008
rect 2626 2944 2643 3008
rect 2707 2944 2724 3008
rect 2788 2944 2805 3008
rect 2869 2944 2886 3008
rect 2950 2944 2967 3008
rect 3031 2944 3048 3008
rect 3112 2944 3129 3008
rect 3193 2944 3210 3008
rect 3274 2944 3291 3008
rect 3355 2944 3372 3008
rect 3436 2944 3453 3008
rect 3517 2944 3534 3008
rect 3598 2944 3615 3008
rect 3679 2944 3696 3008
rect 3760 2944 3777 3008
rect 3841 2944 3858 3008
rect 3922 2944 3939 3008
rect 4003 2944 4020 3008
rect 4084 2944 4101 3008
rect 4165 2944 4182 3008
rect 4246 2944 4263 3008
rect 4327 2944 4344 3008
rect 4408 2944 4425 3008
rect 4489 2944 4506 3008
rect 4570 2944 4587 3008
rect 4651 2944 4668 3008
rect 4732 2944 4749 3008
rect 4813 2944 4830 3008
rect 4894 2944 4895 3008
rect 0 2920 4895 2944
rect 0 2856 126 2920
rect 190 2856 208 2920
rect 272 2856 290 2920
rect 354 2856 372 2920
rect 436 2856 454 2920
rect 518 2856 536 2920
rect 600 2856 618 2920
rect 682 2856 699 2920
rect 763 2856 780 2920
rect 844 2856 861 2920
rect 925 2856 942 2920
rect 1006 2856 1023 2920
rect 1087 2856 1104 2920
rect 1168 2856 1185 2920
rect 1249 2856 1266 2920
rect 1330 2856 1347 2920
rect 1411 2856 1428 2920
rect 1492 2856 1509 2920
rect 1573 2856 1590 2920
rect 1654 2856 1671 2920
rect 1735 2856 1752 2920
rect 1816 2856 1833 2920
rect 1897 2856 1914 2920
rect 1978 2856 1995 2920
rect 2059 2856 2076 2920
rect 2140 2856 2157 2920
rect 2221 2856 2238 2920
rect 2302 2856 2319 2920
rect 2383 2856 2400 2920
rect 2464 2856 2481 2920
rect 2545 2856 2562 2920
rect 2626 2856 2643 2920
rect 2707 2856 2724 2920
rect 2788 2856 2805 2920
rect 2869 2856 2886 2920
rect 2950 2856 2967 2920
rect 3031 2856 3048 2920
rect 3112 2856 3129 2920
rect 3193 2856 3210 2920
rect 3274 2856 3291 2920
rect 3355 2856 3372 2920
rect 3436 2856 3453 2920
rect 3517 2856 3534 2920
rect 3598 2856 3615 2920
rect 3679 2856 3696 2920
rect 3760 2856 3777 2920
rect 3841 2856 3858 2920
rect 3922 2856 3939 2920
rect 4003 2856 4020 2920
rect 4084 2856 4101 2920
rect 4165 2856 4182 2920
rect 4246 2856 4263 2920
rect 4327 2856 4344 2920
rect 4408 2856 4425 2920
rect 4489 2856 4506 2920
rect 4570 2856 4587 2920
rect 4651 2856 4668 2920
rect 4732 2856 4749 2920
rect 4813 2856 4830 2920
rect 4894 2856 4895 2920
rect 0 2832 4895 2856
rect 0 2768 126 2832
rect 190 2768 208 2832
rect 272 2768 290 2832
rect 354 2768 372 2832
rect 436 2768 454 2832
rect 518 2768 536 2832
rect 600 2768 618 2832
rect 682 2768 699 2832
rect 763 2768 780 2832
rect 844 2768 861 2832
rect 925 2768 942 2832
rect 1006 2768 1023 2832
rect 1087 2768 1104 2832
rect 1168 2768 1185 2832
rect 1249 2768 1266 2832
rect 1330 2768 1347 2832
rect 1411 2768 1428 2832
rect 1492 2768 1509 2832
rect 1573 2768 1590 2832
rect 1654 2768 1671 2832
rect 1735 2768 1752 2832
rect 1816 2768 1833 2832
rect 1897 2768 1914 2832
rect 1978 2768 1995 2832
rect 2059 2768 2076 2832
rect 2140 2768 2157 2832
rect 2221 2768 2238 2832
rect 2302 2768 2319 2832
rect 2383 2768 2400 2832
rect 2464 2768 2481 2832
rect 2545 2768 2562 2832
rect 2626 2768 2643 2832
rect 2707 2768 2724 2832
rect 2788 2768 2805 2832
rect 2869 2768 2886 2832
rect 2950 2768 2967 2832
rect 3031 2768 3048 2832
rect 3112 2768 3129 2832
rect 3193 2768 3210 2832
rect 3274 2768 3291 2832
rect 3355 2768 3372 2832
rect 3436 2768 3453 2832
rect 3517 2768 3534 2832
rect 3598 2768 3615 2832
rect 3679 2768 3696 2832
rect 3760 2768 3777 2832
rect 3841 2768 3858 2832
rect 3922 2768 3939 2832
rect 4003 2768 4020 2832
rect 4084 2768 4101 2832
rect 4165 2768 4182 2832
rect 4246 2768 4263 2832
rect 4327 2768 4344 2832
rect 4408 2768 4425 2832
rect 4489 2768 4506 2832
rect 4570 2768 4587 2832
rect 4651 2768 4668 2832
rect 4732 2768 4749 2832
rect 4813 2768 4830 2832
rect 4894 2768 4895 2832
rect 0 2744 4895 2768
rect 0 2680 126 2744
rect 190 2680 208 2744
rect 272 2680 290 2744
rect 354 2680 372 2744
rect 436 2680 454 2744
rect 518 2680 536 2744
rect 600 2680 618 2744
rect 682 2680 699 2744
rect 763 2680 780 2744
rect 844 2680 861 2744
rect 925 2680 942 2744
rect 1006 2680 1023 2744
rect 1087 2680 1104 2744
rect 1168 2680 1185 2744
rect 1249 2680 1266 2744
rect 1330 2680 1347 2744
rect 1411 2680 1428 2744
rect 1492 2680 1509 2744
rect 1573 2680 1590 2744
rect 1654 2680 1671 2744
rect 1735 2680 1752 2744
rect 1816 2680 1833 2744
rect 1897 2680 1914 2744
rect 1978 2680 1995 2744
rect 2059 2680 2076 2744
rect 2140 2680 2157 2744
rect 2221 2680 2238 2744
rect 2302 2680 2319 2744
rect 2383 2680 2400 2744
rect 2464 2680 2481 2744
rect 2545 2680 2562 2744
rect 2626 2680 2643 2744
rect 2707 2680 2724 2744
rect 2788 2680 2805 2744
rect 2869 2680 2886 2744
rect 2950 2680 2967 2744
rect 3031 2680 3048 2744
rect 3112 2680 3129 2744
rect 3193 2680 3210 2744
rect 3274 2680 3291 2744
rect 3355 2680 3372 2744
rect 3436 2680 3453 2744
rect 3517 2680 3534 2744
rect 3598 2680 3615 2744
rect 3679 2680 3696 2744
rect 3760 2680 3777 2744
rect 3841 2680 3858 2744
rect 3922 2680 3939 2744
rect 4003 2680 4020 2744
rect 4084 2680 4101 2744
rect 4165 2680 4182 2744
rect 4246 2680 4263 2744
rect 4327 2680 4344 2744
rect 4408 2680 4425 2744
rect 4489 2680 4506 2744
rect 4570 2680 4587 2744
rect 4651 2680 4668 2744
rect 4732 2680 4749 2744
rect 4813 2680 4830 2744
rect 4894 2680 4895 2744
rect 0 2656 4895 2680
rect 0 2592 126 2656
rect 190 2592 208 2656
rect 272 2592 290 2656
rect 354 2592 372 2656
rect 436 2592 454 2656
rect 518 2592 536 2656
rect 600 2592 618 2656
rect 682 2592 699 2656
rect 763 2592 780 2656
rect 844 2592 861 2656
rect 925 2592 942 2656
rect 1006 2592 1023 2656
rect 1087 2592 1104 2656
rect 1168 2592 1185 2656
rect 1249 2592 1266 2656
rect 1330 2592 1347 2656
rect 1411 2592 1428 2656
rect 1492 2592 1509 2656
rect 1573 2592 1590 2656
rect 1654 2592 1671 2656
rect 1735 2592 1752 2656
rect 1816 2592 1833 2656
rect 1897 2592 1914 2656
rect 1978 2592 1995 2656
rect 2059 2592 2076 2656
rect 2140 2592 2157 2656
rect 2221 2592 2238 2656
rect 2302 2592 2319 2656
rect 2383 2592 2400 2656
rect 2464 2592 2481 2656
rect 2545 2592 2562 2656
rect 2626 2592 2643 2656
rect 2707 2592 2724 2656
rect 2788 2592 2805 2656
rect 2869 2592 2886 2656
rect 2950 2592 2967 2656
rect 3031 2592 3048 2656
rect 3112 2592 3129 2656
rect 3193 2592 3210 2656
rect 3274 2592 3291 2656
rect 3355 2592 3372 2656
rect 3436 2592 3453 2656
rect 3517 2592 3534 2656
rect 3598 2592 3615 2656
rect 3679 2592 3696 2656
rect 3760 2592 3777 2656
rect 3841 2592 3858 2656
rect 3922 2592 3939 2656
rect 4003 2592 4020 2656
rect 4084 2592 4101 2656
rect 4165 2592 4182 2656
rect 4246 2592 4263 2656
rect 4327 2592 4344 2656
rect 4408 2592 4425 2656
rect 4489 2592 4506 2656
rect 4570 2592 4587 2656
rect 4651 2592 4668 2656
rect 4732 2592 4749 2656
rect 4813 2592 4830 2656
rect 4894 2592 4895 2656
rect 0 2587 4895 2592
rect 10156 3272 15000 3277
rect 10156 3208 10157 3272
rect 10221 3208 10239 3272
rect 10303 3208 10321 3272
rect 10385 3208 10403 3272
rect 10467 3208 10485 3272
rect 10549 3208 10567 3272
rect 10631 3208 10649 3272
rect 10713 3208 10730 3272
rect 10794 3208 10811 3272
rect 10875 3208 10892 3272
rect 10956 3208 10973 3272
rect 11037 3208 11054 3272
rect 11118 3208 11135 3272
rect 11199 3208 11216 3272
rect 11280 3208 11297 3272
rect 11361 3208 11378 3272
rect 11442 3208 11459 3272
rect 11523 3208 11540 3272
rect 11604 3208 11621 3272
rect 11685 3208 11702 3272
rect 11766 3208 11783 3272
rect 11847 3208 11864 3272
rect 11928 3208 11945 3272
rect 12009 3208 12026 3272
rect 12090 3208 12107 3272
rect 12171 3208 12188 3272
rect 12252 3208 12269 3272
rect 12333 3208 12350 3272
rect 12414 3208 12431 3272
rect 12495 3208 12512 3272
rect 12576 3208 12593 3272
rect 12657 3208 12674 3272
rect 12738 3208 12755 3272
rect 12819 3208 12836 3272
rect 12900 3208 12917 3272
rect 12981 3208 12998 3272
rect 13062 3208 13079 3272
rect 13143 3208 13160 3272
rect 13224 3208 13241 3272
rect 13305 3208 13322 3272
rect 13386 3208 13403 3272
rect 13467 3208 13484 3272
rect 13548 3208 13565 3272
rect 13629 3208 13646 3272
rect 13710 3208 13727 3272
rect 13791 3208 13808 3272
rect 13872 3208 13889 3272
rect 13953 3208 13970 3272
rect 14034 3208 14051 3272
rect 14115 3208 14132 3272
rect 14196 3208 14213 3272
rect 14277 3208 14294 3272
rect 14358 3208 14375 3272
rect 14439 3208 14456 3272
rect 14520 3208 14537 3272
rect 14601 3208 14618 3272
rect 14682 3208 14699 3272
rect 14763 3208 14780 3272
rect 14844 3208 14861 3272
rect 14925 3208 15000 3272
rect 10156 3184 15000 3208
rect 10156 3120 10157 3184
rect 10221 3120 10239 3184
rect 10303 3120 10321 3184
rect 10385 3120 10403 3184
rect 10467 3120 10485 3184
rect 10549 3120 10567 3184
rect 10631 3120 10649 3184
rect 10713 3120 10730 3184
rect 10794 3120 10811 3184
rect 10875 3120 10892 3184
rect 10956 3120 10973 3184
rect 11037 3120 11054 3184
rect 11118 3120 11135 3184
rect 11199 3120 11216 3184
rect 11280 3120 11297 3184
rect 11361 3120 11378 3184
rect 11442 3120 11459 3184
rect 11523 3120 11540 3184
rect 11604 3120 11621 3184
rect 11685 3120 11702 3184
rect 11766 3120 11783 3184
rect 11847 3120 11864 3184
rect 11928 3120 11945 3184
rect 12009 3120 12026 3184
rect 12090 3120 12107 3184
rect 12171 3120 12188 3184
rect 12252 3120 12269 3184
rect 12333 3120 12350 3184
rect 12414 3120 12431 3184
rect 12495 3120 12512 3184
rect 12576 3120 12593 3184
rect 12657 3120 12674 3184
rect 12738 3120 12755 3184
rect 12819 3120 12836 3184
rect 12900 3120 12917 3184
rect 12981 3120 12998 3184
rect 13062 3120 13079 3184
rect 13143 3120 13160 3184
rect 13224 3120 13241 3184
rect 13305 3120 13322 3184
rect 13386 3120 13403 3184
rect 13467 3120 13484 3184
rect 13548 3120 13565 3184
rect 13629 3120 13646 3184
rect 13710 3120 13727 3184
rect 13791 3120 13808 3184
rect 13872 3120 13889 3184
rect 13953 3120 13970 3184
rect 14034 3120 14051 3184
rect 14115 3120 14132 3184
rect 14196 3120 14213 3184
rect 14277 3120 14294 3184
rect 14358 3120 14375 3184
rect 14439 3120 14456 3184
rect 14520 3120 14537 3184
rect 14601 3120 14618 3184
rect 14682 3120 14699 3184
rect 14763 3120 14780 3184
rect 14844 3120 14861 3184
rect 14925 3120 15000 3184
rect 10156 3096 15000 3120
rect 10156 3032 10157 3096
rect 10221 3032 10239 3096
rect 10303 3032 10321 3096
rect 10385 3032 10403 3096
rect 10467 3032 10485 3096
rect 10549 3032 10567 3096
rect 10631 3032 10649 3096
rect 10713 3032 10730 3096
rect 10794 3032 10811 3096
rect 10875 3032 10892 3096
rect 10956 3032 10973 3096
rect 11037 3032 11054 3096
rect 11118 3032 11135 3096
rect 11199 3032 11216 3096
rect 11280 3032 11297 3096
rect 11361 3032 11378 3096
rect 11442 3032 11459 3096
rect 11523 3032 11540 3096
rect 11604 3032 11621 3096
rect 11685 3032 11702 3096
rect 11766 3032 11783 3096
rect 11847 3032 11864 3096
rect 11928 3032 11945 3096
rect 12009 3032 12026 3096
rect 12090 3032 12107 3096
rect 12171 3032 12188 3096
rect 12252 3032 12269 3096
rect 12333 3032 12350 3096
rect 12414 3032 12431 3096
rect 12495 3032 12512 3096
rect 12576 3032 12593 3096
rect 12657 3032 12674 3096
rect 12738 3032 12755 3096
rect 12819 3032 12836 3096
rect 12900 3032 12917 3096
rect 12981 3032 12998 3096
rect 13062 3032 13079 3096
rect 13143 3032 13160 3096
rect 13224 3032 13241 3096
rect 13305 3032 13322 3096
rect 13386 3032 13403 3096
rect 13467 3032 13484 3096
rect 13548 3032 13565 3096
rect 13629 3032 13646 3096
rect 13710 3032 13727 3096
rect 13791 3032 13808 3096
rect 13872 3032 13889 3096
rect 13953 3032 13970 3096
rect 14034 3032 14051 3096
rect 14115 3032 14132 3096
rect 14196 3032 14213 3096
rect 14277 3032 14294 3096
rect 14358 3032 14375 3096
rect 14439 3032 14456 3096
rect 14520 3032 14537 3096
rect 14601 3032 14618 3096
rect 14682 3032 14699 3096
rect 14763 3032 14780 3096
rect 14844 3032 14861 3096
rect 14925 3032 15000 3096
rect 10156 3008 15000 3032
rect 10156 2944 10157 3008
rect 10221 2944 10239 3008
rect 10303 2944 10321 3008
rect 10385 2944 10403 3008
rect 10467 2944 10485 3008
rect 10549 2944 10567 3008
rect 10631 2944 10649 3008
rect 10713 2944 10730 3008
rect 10794 2944 10811 3008
rect 10875 2944 10892 3008
rect 10956 2944 10973 3008
rect 11037 2944 11054 3008
rect 11118 2944 11135 3008
rect 11199 2944 11216 3008
rect 11280 2944 11297 3008
rect 11361 2944 11378 3008
rect 11442 2944 11459 3008
rect 11523 2944 11540 3008
rect 11604 2944 11621 3008
rect 11685 2944 11702 3008
rect 11766 2944 11783 3008
rect 11847 2944 11864 3008
rect 11928 2944 11945 3008
rect 12009 2944 12026 3008
rect 12090 2944 12107 3008
rect 12171 2944 12188 3008
rect 12252 2944 12269 3008
rect 12333 2944 12350 3008
rect 12414 2944 12431 3008
rect 12495 2944 12512 3008
rect 12576 2944 12593 3008
rect 12657 2944 12674 3008
rect 12738 2944 12755 3008
rect 12819 2944 12836 3008
rect 12900 2944 12917 3008
rect 12981 2944 12998 3008
rect 13062 2944 13079 3008
rect 13143 2944 13160 3008
rect 13224 2944 13241 3008
rect 13305 2944 13322 3008
rect 13386 2944 13403 3008
rect 13467 2944 13484 3008
rect 13548 2944 13565 3008
rect 13629 2944 13646 3008
rect 13710 2944 13727 3008
rect 13791 2944 13808 3008
rect 13872 2944 13889 3008
rect 13953 2944 13970 3008
rect 14034 2944 14051 3008
rect 14115 2944 14132 3008
rect 14196 2944 14213 3008
rect 14277 2944 14294 3008
rect 14358 2944 14375 3008
rect 14439 2944 14456 3008
rect 14520 2944 14537 3008
rect 14601 2944 14618 3008
rect 14682 2944 14699 3008
rect 14763 2944 14780 3008
rect 14844 2944 14861 3008
rect 14925 2944 15000 3008
rect 10156 2920 15000 2944
rect 10156 2856 10157 2920
rect 10221 2856 10239 2920
rect 10303 2856 10321 2920
rect 10385 2856 10403 2920
rect 10467 2856 10485 2920
rect 10549 2856 10567 2920
rect 10631 2856 10649 2920
rect 10713 2856 10730 2920
rect 10794 2856 10811 2920
rect 10875 2856 10892 2920
rect 10956 2856 10973 2920
rect 11037 2856 11054 2920
rect 11118 2856 11135 2920
rect 11199 2856 11216 2920
rect 11280 2856 11297 2920
rect 11361 2856 11378 2920
rect 11442 2856 11459 2920
rect 11523 2856 11540 2920
rect 11604 2856 11621 2920
rect 11685 2856 11702 2920
rect 11766 2856 11783 2920
rect 11847 2856 11864 2920
rect 11928 2856 11945 2920
rect 12009 2856 12026 2920
rect 12090 2856 12107 2920
rect 12171 2856 12188 2920
rect 12252 2856 12269 2920
rect 12333 2856 12350 2920
rect 12414 2856 12431 2920
rect 12495 2856 12512 2920
rect 12576 2856 12593 2920
rect 12657 2856 12674 2920
rect 12738 2856 12755 2920
rect 12819 2856 12836 2920
rect 12900 2856 12917 2920
rect 12981 2856 12998 2920
rect 13062 2856 13079 2920
rect 13143 2856 13160 2920
rect 13224 2856 13241 2920
rect 13305 2856 13322 2920
rect 13386 2856 13403 2920
rect 13467 2856 13484 2920
rect 13548 2856 13565 2920
rect 13629 2856 13646 2920
rect 13710 2856 13727 2920
rect 13791 2856 13808 2920
rect 13872 2856 13889 2920
rect 13953 2856 13970 2920
rect 14034 2856 14051 2920
rect 14115 2856 14132 2920
rect 14196 2856 14213 2920
rect 14277 2856 14294 2920
rect 14358 2856 14375 2920
rect 14439 2856 14456 2920
rect 14520 2856 14537 2920
rect 14601 2856 14618 2920
rect 14682 2856 14699 2920
rect 14763 2856 14780 2920
rect 14844 2856 14861 2920
rect 14925 2856 15000 2920
rect 10156 2832 15000 2856
rect 10156 2768 10157 2832
rect 10221 2768 10239 2832
rect 10303 2768 10321 2832
rect 10385 2768 10403 2832
rect 10467 2768 10485 2832
rect 10549 2768 10567 2832
rect 10631 2768 10649 2832
rect 10713 2768 10730 2832
rect 10794 2768 10811 2832
rect 10875 2768 10892 2832
rect 10956 2768 10973 2832
rect 11037 2768 11054 2832
rect 11118 2768 11135 2832
rect 11199 2768 11216 2832
rect 11280 2768 11297 2832
rect 11361 2768 11378 2832
rect 11442 2768 11459 2832
rect 11523 2768 11540 2832
rect 11604 2768 11621 2832
rect 11685 2768 11702 2832
rect 11766 2768 11783 2832
rect 11847 2768 11864 2832
rect 11928 2768 11945 2832
rect 12009 2768 12026 2832
rect 12090 2768 12107 2832
rect 12171 2768 12188 2832
rect 12252 2768 12269 2832
rect 12333 2768 12350 2832
rect 12414 2768 12431 2832
rect 12495 2768 12512 2832
rect 12576 2768 12593 2832
rect 12657 2768 12674 2832
rect 12738 2768 12755 2832
rect 12819 2768 12836 2832
rect 12900 2768 12917 2832
rect 12981 2768 12998 2832
rect 13062 2768 13079 2832
rect 13143 2768 13160 2832
rect 13224 2768 13241 2832
rect 13305 2768 13322 2832
rect 13386 2768 13403 2832
rect 13467 2768 13484 2832
rect 13548 2768 13565 2832
rect 13629 2768 13646 2832
rect 13710 2768 13727 2832
rect 13791 2768 13808 2832
rect 13872 2768 13889 2832
rect 13953 2768 13970 2832
rect 14034 2768 14051 2832
rect 14115 2768 14132 2832
rect 14196 2768 14213 2832
rect 14277 2768 14294 2832
rect 14358 2768 14375 2832
rect 14439 2768 14456 2832
rect 14520 2768 14537 2832
rect 14601 2768 14618 2832
rect 14682 2768 14699 2832
rect 14763 2768 14780 2832
rect 14844 2768 14861 2832
rect 14925 2768 15000 2832
rect 10156 2744 15000 2768
rect 10156 2680 10157 2744
rect 10221 2680 10239 2744
rect 10303 2680 10321 2744
rect 10385 2680 10403 2744
rect 10467 2680 10485 2744
rect 10549 2680 10567 2744
rect 10631 2680 10649 2744
rect 10713 2680 10730 2744
rect 10794 2680 10811 2744
rect 10875 2680 10892 2744
rect 10956 2680 10973 2744
rect 11037 2680 11054 2744
rect 11118 2680 11135 2744
rect 11199 2680 11216 2744
rect 11280 2680 11297 2744
rect 11361 2680 11378 2744
rect 11442 2680 11459 2744
rect 11523 2680 11540 2744
rect 11604 2680 11621 2744
rect 11685 2680 11702 2744
rect 11766 2680 11783 2744
rect 11847 2680 11864 2744
rect 11928 2680 11945 2744
rect 12009 2680 12026 2744
rect 12090 2680 12107 2744
rect 12171 2680 12188 2744
rect 12252 2680 12269 2744
rect 12333 2680 12350 2744
rect 12414 2680 12431 2744
rect 12495 2680 12512 2744
rect 12576 2680 12593 2744
rect 12657 2680 12674 2744
rect 12738 2680 12755 2744
rect 12819 2680 12836 2744
rect 12900 2680 12917 2744
rect 12981 2680 12998 2744
rect 13062 2680 13079 2744
rect 13143 2680 13160 2744
rect 13224 2680 13241 2744
rect 13305 2680 13322 2744
rect 13386 2680 13403 2744
rect 13467 2680 13484 2744
rect 13548 2680 13565 2744
rect 13629 2680 13646 2744
rect 13710 2680 13727 2744
rect 13791 2680 13808 2744
rect 13872 2680 13889 2744
rect 13953 2680 13970 2744
rect 14034 2680 14051 2744
rect 14115 2680 14132 2744
rect 14196 2680 14213 2744
rect 14277 2680 14294 2744
rect 14358 2680 14375 2744
rect 14439 2680 14456 2744
rect 14520 2680 14537 2744
rect 14601 2680 14618 2744
rect 14682 2680 14699 2744
rect 14763 2680 14780 2744
rect 14844 2680 14861 2744
rect 14925 2680 15000 2744
rect 10156 2656 15000 2680
rect 10156 2592 10157 2656
rect 10221 2592 10239 2656
rect 10303 2592 10321 2656
rect 10385 2592 10403 2656
rect 10467 2592 10485 2656
rect 10549 2592 10567 2656
rect 10631 2592 10649 2656
rect 10713 2592 10730 2656
rect 10794 2592 10811 2656
rect 10875 2592 10892 2656
rect 10956 2592 10973 2656
rect 11037 2592 11054 2656
rect 11118 2592 11135 2656
rect 11199 2592 11216 2656
rect 11280 2592 11297 2656
rect 11361 2592 11378 2656
rect 11442 2592 11459 2656
rect 11523 2592 11540 2656
rect 11604 2592 11621 2656
rect 11685 2592 11702 2656
rect 11766 2592 11783 2656
rect 11847 2592 11864 2656
rect 11928 2592 11945 2656
rect 12009 2592 12026 2656
rect 12090 2592 12107 2656
rect 12171 2592 12188 2656
rect 12252 2592 12269 2656
rect 12333 2592 12350 2656
rect 12414 2592 12431 2656
rect 12495 2592 12512 2656
rect 12576 2592 12593 2656
rect 12657 2592 12674 2656
rect 12738 2592 12755 2656
rect 12819 2592 12836 2656
rect 12900 2592 12917 2656
rect 12981 2592 12998 2656
rect 13062 2592 13079 2656
rect 13143 2592 13160 2656
rect 13224 2592 13241 2656
rect 13305 2592 13322 2656
rect 13386 2592 13403 2656
rect 13467 2592 13484 2656
rect 13548 2592 13565 2656
rect 13629 2592 13646 2656
rect 13710 2592 13727 2656
rect 13791 2592 13808 2656
rect 13872 2592 13889 2656
rect 13953 2592 13970 2656
rect 14034 2592 14051 2656
rect 14115 2592 14132 2656
rect 14196 2592 14213 2656
rect 14277 2592 14294 2656
rect 14358 2592 14375 2656
rect 14439 2592 14456 2656
rect 14520 2592 14537 2656
rect 14601 2592 14618 2656
rect 14682 2592 14699 2656
rect 14763 2592 14780 2656
rect 14844 2592 14861 2656
rect 14925 2592 15000 2656
rect 10156 2587 15000 2592
rect 0 1377 254 2307
rect 14746 1377 15000 2307
rect 0 7 254 1097
rect 14746 7 15000 1097
<< metal5 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18597
rect 14746 13607 15000 18597
rect 0 12437 254 13287
rect 14746 12437 15000 13287
rect 0 11267 254 12117
rect 14746 11267 15000 12117
rect 0 9147 254 10947
rect 14746 9147 15000 10947
rect 0 7937 254 8827
rect 14746 7937 15000 8827
rect 0 6968 254 7617
rect 14746 6968 15000 7617
rect 0 5997 254 6647
rect 14746 5997 15000 6647
rect 0 4787 254 5677
rect 14746 4787 15000 5677
rect 0 3577 254 4467
rect 14746 3577 15000 4467
rect 0 2607 193 3257
rect 14807 2607 15000 3257
rect 0 1397 254 2287
rect 14746 1397 15000 2287
rect 0 27 254 1077
rect 14746 27 15000 1077
use sky130_fd_io__com_bus_hookup  sky130_fd_io__com_bus_hookup_0
timestamp 1683767628
transform 1 0 0 0 1 149
box 0 -142 15000 39451
<< labels >>
flabel metal5 s 0 5997 254 6647 3 FreeSans 520 0 0 0 VSWITCH
port 1 nsew power bidirectional
flabel metal5 s 14746 5997 15000 6647 3 FreeSans 520 180 0 0 VSWITCH
port 1 nsew power bidirectional
flabel metal5 s 0 1397 254 2287 3 FreeSans 520 0 0 0 VCCD
port 2 nsew power bidirectional
flabel metal5 s 0 27 254 1077 3 FreeSans 520 0 0 0 VCCHIB
port 3 nsew power bidirectional
flabel metal5 s 14807 2607 15000 3257 3 FreeSans 520 180 0 0 VDDA
port 4 nsew power bidirectional
flabel metal5 s 0 2607 193 3257 3 FreeSans 520 0 0 0 VDDA
port 4 nsew power bidirectional
flabel metal5 s 14746 7937 15000 8827 3 FreeSans 520 180 0 0 VSSD
port 5 nsew ground bidirectional
flabel metal5 s 14746 13607 15000 18597 3 FreeSans 520 180 0 0 VDDIO
port 6 nsew power bidirectional
flabel metal5 s 0 13607 254 18597 3 FreeSans 520 0 0 0 VDDIO
port 6 nsew power bidirectional
flabel metal5 s 0 3577 254 4467 3 FreeSans 520 0 0 0 VDDIO
port 6 nsew power bidirectional
flabel metal5 s 14746 12437 15000 13287 3 FreeSans 520 180 0 0 VDDIO_Q
port 7 nsew power bidirectional
flabel metal5 s 14746 9147 15000 10947 3 FreeSans 520 180 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal5 s 14746 6968 15000 7617 3 FreeSans 520 180 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal5 s 0 9147 254 10947 3 FreeSans 520 0 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal5 s 0 6968 254 7617 3 FreeSans 520 0 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal5 s 0 7937 254 8827 3 FreeSans 520 0 0 0 VSSD
port 5 nsew ground bidirectional
flabel metal5 s 14746 34757 15000 39600 3 FreeSans 520 180 0 0 VSSIO
port 9 nsew ground bidirectional
flabel metal5 s 0 12437 254 13287 3 FreeSans 520 0 0 0 VDDIO_Q
port 7 nsew power bidirectional
flabel metal5 s 14746 4787 15000 5677 3 FreeSans 520 180 0 0 VSSIO
port 9 nsew ground bidirectional
flabel metal5 s 14746 1397 15000 2287 3 FreeSans 520 180 0 0 VCCD
port 2 nsew power bidirectional
flabel metal5 s 14746 27 15000 1077 3 FreeSans 520 180 0 0 VCCHIB
port 3 nsew power bidirectional
flabel metal5 s 0 34757 254 39600 3 FreeSans 520 0 0 0 VSSIO
port 9 nsew ground bidirectional
flabel metal5 s 14746 3577 15000 4467 3 FreeSans 520 180 0 0 VDDIO
port 6 nsew power bidirectional
flabel metal5 s 0 4787 254 5677 3 FreeSans 520 0 0 0 VSSIO
port 9 nsew ground bidirectional
flabel metal5 s 14746 11267 15000 12117 3 FreeSans 520 180 0 0 VSSIO_Q
port 10 nsew ground bidirectional
flabel metal5 s 0 11267 254 12117 3 FreeSans 520 0 0 0 VSSIO_Q
port 10 nsew ground bidirectional
flabel metal4 s 0 5977 254 6667 3 FreeSans 520 0 0 0 VSWITCH
port 1 nsew power bidirectional
flabel metal4 s 14746 5977 15000 6667 3 FreeSans 520 180 0 0 VSWITCH
port 1 nsew power bidirectional
flabel metal4 s 14746 10225 15000 10821 3 FreeSans 520 180 0 0 AMUXBUS_A
port 12 nsew signal bidirectional
flabel metal4 s 0 10225 254 10821 3 FreeSans 520 0 0 0 AMUXBUS_A
port 12 nsew signal bidirectional
flabel metal4 s 14746 9273 15000 9869 3 FreeSans 520 180 0 0 AMUXBUS_B
port 11 nsew signal bidirectional
flabel metal4 s 14746 1377 15000 2307 3 FreeSans 520 180 0 0 VCCD
port 2 nsew power bidirectional
flabel metal4 s 0 1377 254 2307 3 FreeSans 520 0 0 0 VCCD
port 2 nsew power bidirectional
flabel metal4 s 14746 7 15000 1097 3 FreeSans 520 180 0 0 VCCHIB
port 3 nsew power bidirectional
flabel metal4 s 0 7 254 1097 3 FreeSans 520 0 0 0 VCCHIB
port 3 nsew power bidirectional
flabel metal4 s 14807 2587 15000 3277 3 FreeSans 520 180 0 0 VDDA
port 4 nsew power bidirectional
flabel metal4 s 0 2587 193 3277 3 FreeSans 520 0 0 0 VDDA
port 4 nsew power bidirectional
flabel metal4 s 14746 3557 15000 4487 3 FreeSans 520 180 0 0 VDDIO
port 6 nsew power bidirectional
flabel metal4 s 14746 7917 15000 8847 3 FreeSans 520 180 0 0 VSSD
port 5 nsew ground bidirectional
flabel metal4 s 14746 13607 15000 18600 3 FreeSans 520 180 0 0 VDDIO
port 6 nsew power bidirectional
flabel metal4 s 0 3557 254 4487 3 FreeSans 520 0 0 0 VDDIO
port 6 nsew power bidirectional
flabel metal4 s 0 13607 254 18600 3 FreeSans 520 0 0 0 VDDIO
port 6 nsew power bidirectional
flabel metal4 s 14746 12417 15000 13307 3 FreeSans 520 180 0 0 VDDIO_Q
port 7 nsew power bidirectional
flabel metal4 s 14746 6947 15000 7637 3 FreeSans 520 180 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal4 s 14746 9147 15000 9213 3 FreeSans 520 180 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal4 s 14746 10881 15000 10947 3 FreeSans 520 180 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal4 s 14746 9929 15000 10165 3 FreeSans 520 180 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal4 s 0 9147 254 9213 3 FreeSans 520 0 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal4 s 0 9929 254 10165 3 FreeSans 520 0 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal4 s 0 10881 254 10947 3 FreeSans 520 0 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal4 s 0 6947 254 7637 3 FreeSans 520 0 0 0 VSSA
port 8 nsew ground bidirectional
flabel metal4 s 0 7917 254 8847 3 FreeSans 520 0 0 0 VSSD
port 5 nsew ground bidirectional
flabel metal4 s 14746 34757 15000 39600 3 FreeSans 520 180 0 0 VSSIO
port 9 nsew ground bidirectional
flabel metal4 s 0 9273 254 9869 3 FreeSans 520 0 0 0 AMUXBUS_B
port 11 nsew signal bidirectional
flabel metal4 s 14746 4767 15000 5697 3 FreeSans 520 180 0 0 VSSIO
port 9 nsew ground bidirectional
flabel metal4 s 0 12417 254 13307 3 FreeSans 520 0 0 0 VDDIO_Q
port 7 nsew power bidirectional
flabel metal4 s 0 34757 254 39600 3 FreeSans 520 0 0 0 VSSIO
port 9 nsew ground bidirectional
flabel metal4 s 0 4767 254 5697 3 FreeSans 520 0 0 0 VSSIO
port 9 nsew ground bidirectional
flabel metal4 s 14746 11247 15000 12137 3 FreeSans 520 180 0 0 VSSIO_Q
port 10 nsew ground bidirectional
flabel metal4 s 0 11247 254 12137 3 FreeSans 520 0 0 0 VSSIO_Q
port 10 nsew ground bidirectional
rlabel metal4 s 14746 10225 15000 10821 1 AMUXBUS_A
port 12 nsew signal bidirectional
rlabel metal4 s 14746 9273 15000 9869 1 AMUXBUS_B
port 11 nsew signal bidirectional
rlabel metal4 s 14746 1377 15000 2307 1 VCCD
port 2 nsew power bidirectional
rlabel metal5 s 0 1397 254 2287 1 VCCD
port 2 nsew power bidirectional
rlabel metal5 s 14746 1397 15000 2287 1 VCCD
port 2 nsew power bidirectional
rlabel metal4 s 14746 7 15000 1097 1 VCCHIB
port 3 nsew power bidirectional
rlabel metal5 s 0 27 254 1077 1 VCCHIB
port 3 nsew power bidirectional
rlabel metal5 s 14746 27 15000 1077 1 VCCHIB
port 3 nsew power bidirectional
rlabel metal3 s 10151 2588 14931 3276 1 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 0 2587 4895 3277 1 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 10156 2587 15000 3277 1 VDDA
port 4 nsew power bidirectional
rlabel metal5 s 0 2607 193 3257 1 VDDA
port 4 nsew power bidirectional
rlabel metal5 s 14807 2607 15000 3257 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14873 3220 14913 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14873 3132 14913 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14873 3044 14913 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14873 2956 14913 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14873 2868 14913 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14873 2780 14913 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14873 2692 14913 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14873 2604 14913 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14792 3220 14832 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14792 3132 14832 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14792 3044 14832 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14792 2956 14832 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14792 2868 14832 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14792 2780 14832 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14792 2692 14832 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14792 2604 14832 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14711 3220 14751 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14711 3132 14751 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14711 3044 14751 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14711 2956 14751 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14711 2868 14751 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14711 2780 14751 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14711 2692 14751 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14711 2604 14751 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14630 3220 14670 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14630 3132 14670 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14630 3044 14670 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14630 2956 14670 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14630 2868 14670 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14630 2780 14670 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14630 2692 14670 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14630 2604 14670 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14549 3220 14589 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14549 3132 14589 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14549 3044 14589 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14549 2956 14589 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14549 2868 14589 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14549 2780 14589 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14549 2692 14589 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14549 2604 14589 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14468 3220 14508 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14468 3132 14508 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14468 3044 14508 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14468 2956 14508 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14468 2868 14508 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14468 2780 14508 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14468 2692 14508 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14468 2604 14508 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14387 3220 14427 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14387 3132 14427 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14387 3044 14427 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14387 2956 14427 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14387 2868 14427 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14387 2780 14427 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14387 2692 14427 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14387 2604 14427 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14306 3220 14346 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14306 3132 14346 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14306 3044 14346 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14306 2956 14346 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14306 2868 14346 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14306 2780 14346 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14306 2692 14346 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14306 2604 14346 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14225 3220 14265 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14225 3132 14265 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14225 3044 14265 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14225 2956 14265 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14225 2868 14265 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14225 2780 14265 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14225 2692 14265 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14225 2604 14265 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14144 3220 14184 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14144 3132 14184 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14144 3044 14184 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14144 2956 14184 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14144 2868 14184 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14144 2780 14184 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14144 2692 14184 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14144 2604 14184 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14063 3220 14103 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14063 3132 14103 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14063 3044 14103 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14063 2956 14103 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14063 2868 14103 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14063 2780 14103 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14063 2692 14103 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 14063 2604 14103 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13982 3220 14022 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13982 3132 14022 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13982 3044 14022 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13982 2956 14022 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13982 2868 14022 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13982 2780 14022 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13982 2692 14022 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13982 2604 14022 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13901 3220 13941 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13901 3132 13941 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13901 3044 13941 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13901 2956 13941 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13901 2868 13941 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13901 2780 13941 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13901 2692 13941 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13901 2604 13941 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13820 3220 13860 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13820 3132 13860 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13820 3044 13860 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13820 2956 13860 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13820 2868 13860 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13820 2780 13860 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13820 2692 13860 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13820 2604 13860 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13739 3220 13779 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13739 3132 13779 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13739 3044 13779 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13739 2956 13779 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13739 2868 13779 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13739 2780 13779 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13739 2692 13779 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13739 2604 13779 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13658 3220 13698 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13658 3132 13698 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13658 3044 13698 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13658 2956 13698 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13658 2868 13698 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13658 2780 13698 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13658 2692 13698 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13658 2604 13698 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13577 3220 13617 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13577 3132 13617 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13577 3044 13617 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13577 2956 13617 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13577 2868 13617 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13577 2780 13617 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13577 2692 13617 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13577 2604 13617 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13496 3220 13536 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13496 3132 13536 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13496 3044 13536 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13496 2956 13536 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13496 2868 13536 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13496 2780 13536 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13496 2692 13536 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13496 2604 13536 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13415 3220 13455 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13415 3132 13455 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13415 3044 13455 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13415 2956 13455 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13415 2868 13455 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13415 2780 13455 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13415 2692 13455 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13415 2604 13455 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13334 3220 13374 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13334 3132 13374 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13334 3044 13374 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13334 2956 13374 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13334 2868 13374 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13334 2780 13374 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13334 2692 13374 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13334 2604 13374 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13253 3220 13293 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13253 3132 13293 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13253 3044 13293 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13253 2956 13293 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13253 2868 13293 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13253 2780 13293 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13253 2692 13293 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13253 2604 13293 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13172 3220 13212 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13172 3132 13212 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13172 3044 13212 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13172 2956 13212 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13172 2868 13212 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13172 2780 13212 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13172 2692 13212 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13172 2604 13212 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13091 3220 13131 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13091 3132 13131 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13091 3044 13131 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13091 2956 13131 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13091 2868 13131 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13091 2780 13131 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13091 2692 13131 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13091 2604 13131 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13010 3220 13050 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13010 3132 13050 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13010 3044 13050 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13010 2956 13050 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13010 2868 13050 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13010 2780 13050 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13010 2692 13050 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 13010 2604 13050 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12929 3220 12969 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12929 3132 12969 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12929 3044 12969 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12929 2956 12969 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12929 2868 12969 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12929 2780 12969 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12929 2692 12969 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12929 2604 12969 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12848 3220 12888 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12848 3132 12888 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12848 3044 12888 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12848 2956 12888 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12848 2868 12888 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12848 2780 12888 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12848 2692 12888 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12848 2604 12888 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12767 3220 12807 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12767 3132 12807 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12767 3044 12807 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12767 2956 12807 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12767 2868 12807 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12767 2780 12807 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12767 2692 12807 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12767 2604 12807 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12686 3220 12726 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12686 3132 12726 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12686 3044 12726 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12686 2956 12726 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12686 2868 12726 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12686 2780 12726 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12686 2692 12726 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12686 2604 12726 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12605 3220 12645 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12605 3132 12645 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12605 3044 12645 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12605 2956 12645 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12605 2868 12645 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12605 2780 12645 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12605 2692 12645 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12605 2604 12645 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12524 3220 12564 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12524 3132 12564 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12524 3044 12564 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12524 2956 12564 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12524 2868 12564 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12524 2780 12564 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12524 2692 12564 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12524 2604 12564 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12443 3220 12483 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12443 3132 12483 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12443 3044 12483 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12443 2956 12483 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12443 2868 12483 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12443 2780 12483 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12443 2692 12483 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12443 2604 12483 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12362 3220 12402 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12362 3132 12402 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12362 3044 12402 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12362 2956 12402 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12362 2868 12402 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12362 2780 12402 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12362 2692 12402 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12362 2604 12402 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12281 3220 12321 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12281 3132 12321 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12281 3044 12321 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12281 2956 12321 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12281 2868 12321 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12281 2780 12321 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12281 2692 12321 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12281 2604 12321 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12200 3220 12240 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12200 3132 12240 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12200 3044 12240 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12200 2956 12240 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12200 2868 12240 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12200 2780 12240 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12200 2692 12240 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12200 2604 12240 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12119 3220 12159 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12119 3132 12159 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12119 3044 12159 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12119 2956 12159 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12119 2868 12159 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12119 2780 12159 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12119 2692 12159 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12119 2604 12159 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12038 3220 12078 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12038 3132 12078 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12038 3044 12078 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12038 2956 12078 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12038 2868 12078 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12038 2780 12078 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12038 2692 12078 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 12038 2604 12078 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11957 3220 11997 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11957 3132 11997 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11957 3044 11997 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11957 2956 11997 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11957 2868 11997 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11957 2780 11997 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11957 2692 11997 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11957 2604 11997 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11876 3220 11916 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11876 3132 11916 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11876 3044 11916 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11876 2956 11916 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11876 2868 11916 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11876 2780 11916 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11876 2692 11916 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11876 2604 11916 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11795 3220 11835 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11795 3132 11835 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11795 3044 11835 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11795 2956 11835 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11795 2868 11835 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11795 2780 11835 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11795 2692 11835 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11795 2604 11835 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11714 3220 11754 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11714 3132 11754 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11714 3044 11754 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11714 2956 11754 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11714 2868 11754 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11714 2780 11754 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11714 2692 11754 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11714 2604 11754 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11633 3220 11673 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11633 3132 11673 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11633 3044 11673 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11633 2956 11673 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11633 2868 11673 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11633 2780 11673 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11633 2692 11673 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11633 2604 11673 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11552 3220 11592 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11552 3132 11592 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11552 3044 11592 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11552 2956 11592 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11552 2868 11592 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11552 2780 11592 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11552 2692 11592 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11552 2604 11592 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11471 3220 11511 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11471 3132 11511 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11471 3044 11511 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11471 2956 11511 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11471 2868 11511 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11471 2780 11511 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11471 2692 11511 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11471 2604 11511 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11390 3220 11430 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11390 3132 11430 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11390 3044 11430 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11390 2956 11430 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11390 2868 11430 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11390 2780 11430 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11390 2692 11430 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11390 2604 11430 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11309 3220 11349 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11309 3132 11349 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11309 3044 11349 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11309 2956 11349 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11309 2868 11349 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11309 2780 11349 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11309 2692 11349 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11309 2604 11349 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11228 3220 11268 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11228 3132 11268 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11228 3044 11268 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11228 2956 11268 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11228 2868 11268 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11228 2780 11268 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11228 2692 11268 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11228 2604 11268 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11147 3220 11187 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11147 3132 11187 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11147 3044 11187 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11147 2956 11187 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11147 2868 11187 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11147 2780 11187 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11147 2692 11187 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11147 2604 11187 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11066 3220 11106 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11066 3132 11106 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11066 3044 11106 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11066 2956 11106 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11066 2868 11106 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11066 2780 11106 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11066 2692 11106 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 11066 2604 11106 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10985 3220 11025 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10985 3132 11025 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10985 3044 11025 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10985 2956 11025 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10985 2868 11025 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10985 2780 11025 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10985 2692 11025 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10985 2604 11025 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10904 3220 10944 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10904 3132 10944 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10904 3044 10944 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10904 2956 10944 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10904 2868 10944 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10904 2780 10944 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10904 2692 10944 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10904 2604 10944 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10823 3220 10863 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10823 3132 10863 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10823 3044 10863 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10823 2956 10863 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10823 2868 10863 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10823 2780 10863 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10823 2692 10863 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10823 2604 10863 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10742 3220 10782 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10742 3132 10782 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10742 3044 10782 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10742 2956 10782 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10742 2868 10782 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10742 2780 10782 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10742 2692 10782 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10742 2604 10782 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10661 3220 10701 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10661 3132 10701 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10661 3044 10701 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10661 2956 10701 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10661 2868 10701 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10661 2780 10701 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10661 2692 10701 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10661 2604 10701 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10579 3220 10619 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10579 3132 10619 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10579 3044 10619 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10579 2956 10619 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10579 2868 10619 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10579 2780 10619 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10579 2692 10619 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10579 2604 10619 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10497 3220 10537 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10497 3132 10537 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10497 3044 10537 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10497 2956 10537 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10497 2868 10537 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10497 2780 10537 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10497 2692 10537 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10497 2604 10537 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10415 3220 10455 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10415 3132 10455 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10415 3044 10455 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10415 2956 10455 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10415 2868 10455 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10415 2780 10455 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10415 2692 10455 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10415 2604 10455 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10333 3220 10373 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10333 3132 10373 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10333 3044 10373 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10333 2956 10373 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10333 2868 10373 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10333 2780 10373 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10333 2692 10373 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10333 2604 10373 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10251 3220 10291 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10251 3132 10291 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10251 3044 10291 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10251 2956 10291 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10251 2868 10291 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10251 2780 10291 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10251 2692 10291 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10251 2604 10291 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10169 3220 10209 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10169 3132 10209 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10169 3044 10209 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10169 2956 10209 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10169 2868 10209 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10169 2780 10209 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10169 2692 10209 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 10169 2604 10209 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4842 3220 4882 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4842 3132 4882 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4842 3044 4882 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4842 2956 4882 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4842 2868 4882 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4842 2780 4882 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4842 2692 4882 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4842 2604 4882 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4761 3220 4801 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4761 3132 4801 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4761 3044 4801 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4761 2956 4801 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4761 2868 4801 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4761 2780 4801 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4761 2692 4801 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4761 2604 4801 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4680 3220 4720 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4680 3132 4720 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4680 3044 4720 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4680 2956 4720 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4680 2868 4720 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4680 2780 4720 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4680 2692 4720 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4680 2604 4720 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4599 3220 4639 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4599 3132 4639 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4599 3044 4639 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4599 2956 4639 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4599 2868 4639 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4599 2780 4639 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4599 2692 4639 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4599 2604 4639 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4518 3220 4558 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4518 3132 4558 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4518 3044 4558 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4518 2956 4558 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4518 2868 4558 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4518 2780 4558 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4518 2692 4558 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4518 2604 4558 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4437 3220 4477 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4437 3132 4477 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4437 3044 4477 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4437 2956 4477 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4437 2868 4477 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4437 2780 4477 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4437 2692 4477 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4437 2604 4477 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4356 3220 4396 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4356 3132 4396 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4356 3044 4396 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4356 2956 4396 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4356 2868 4396 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4356 2780 4396 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4356 2692 4396 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4356 2604 4396 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4275 3220 4315 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4275 3132 4315 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4275 3044 4315 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4275 2956 4315 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4275 2868 4315 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4275 2780 4315 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4275 2692 4315 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4275 2604 4315 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4194 3220 4234 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4194 3132 4234 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4194 3044 4234 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4194 2956 4234 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4194 2868 4234 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4194 2780 4234 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4194 2692 4234 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4194 2604 4234 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4113 3220 4153 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4113 3132 4153 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4113 3044 4153 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4113 2956 4153 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4113 2868 4153 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4113 2780 4153 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4113 2692 4153 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4113 2604 4153 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4032 3220 4072 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4032 3132 4072 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4032 3044 4072 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4032 2956 4072 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4032 2868 4072 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4032 2780 4072 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4032 2692 4072 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 4032 2604 4072 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3951 3220 3991 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3951 3132 3991 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3951 3044 3991 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3951 2956 3991 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3951 2868 3991 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3951 2780 3991 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3951 2692 3991 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3951 2604 3991 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3870 3220 3910 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3870 3132 3910 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3870 3044 3910 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3870 2956 3910 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3870 2868 3910 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3870 2780 3910 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3870 2692 3910 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3870 2604 3910 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3789 3220 3829 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3789 3132 3829 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3789 3044 3829 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3789 2956 3829 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3789 2868 3829 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3789 2780 3829 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3789 2692 3829 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3789 2604 3829 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3708 3220 3748 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3708 3132 3748 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3708 3044 3748 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3708 2956 3748 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3708 2868 3748 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3708 2780 3748 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3708 2692 3748 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3708 2604 3748 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3627 3220 3667 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3627 3132 3667 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3627 3044 3667 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3627 2956 3667 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3627 2868 3667 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3627 2780 3667 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3627 2692 3667 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3627 2604 3667 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3546 3220 3586 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3546 3132 3586 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3546 3044 3586 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3546 2956 3586 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3546 2868 3586 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3546 2780 3586 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3546 2692 3586 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3546 2604 3586 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3465 3220 3505 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3465 3132 3505 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3465 3044 3505 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3465 2956 3505 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3465 2868 3505 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3465 2780 3505 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3465 2692 3505 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3465 2604 3505 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3384 3220 3424 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3384 3132 3424 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3384 3044 3424 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3384 2956 3424 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3384 2868 3424 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3384 2780 3424 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3384 2692 3424 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3384 2604 3424 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3303 3220 3343 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3303 3132 3343 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3303 3044 3343 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3303 2956 3343 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3303 2868 3343 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3303 2780 3343 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3303 2692 3343 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3303 2604 3343 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3222 3220 3262 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3222 3132 3262 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3222 3044 3262 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3222 2956 3262 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3222 2868 3262 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3222 2780 3262 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3222 2692 3262 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3222 2604 3262 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3141 3220 3181 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3141 3132 3181 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3141 3044 3181 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3141 2956 3181 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3141 2868 3181 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3141 2780 3181 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3141 2692 3181 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3141 2604 3181 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3060 3220 3100 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3060 3132 3100 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3060 3044 3100 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3060 2956 3100 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3060 2868 3100 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3060 2780 3100 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3060 2692 3100 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 3060 2604 3100 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2979 3220 3019 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2979 3132 3019 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2979 3044 3019 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2979 2956 3019 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2979 2868 3019 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2979 2780 3019 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2979 2692 3019 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2979 2604 3019 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2898 3220 2938 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2898 3132 2938 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2898 3044 2938 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2898 2956 2938 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2898 2868 2938 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2898 2780 2938 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2898 2692 2938 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2898 2604 2938 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2817 3220 2857 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2817 3132 2857 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2817 3044 2857 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2817 2956 2857 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2817 2868 2857 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2817 2780 2857 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2817 2692 2857 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2817 2604 2857 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2736 3220 2776 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2736 3132 2776 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2736 3044 2776 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2736 2956 2776 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2736 2868 2776 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2736 2780 2776 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2736 2692 2776 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2736 2604 2776 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2655 3220 2695 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2655 3132 2695 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2655 3044 2695 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2655 2956 2695 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2655 2868 2695 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2655 2780 2695 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2655 2692 2695 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2655 2604 2695 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2574 3220 2614 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2574 3132 2614 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2574 3044 2614 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2574 2956 2614 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2574 2868 2614 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2574 2780 2614 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2574 2692 2614 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2574 2604 2614 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2493 3220 2533 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2493 3132 2533 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2493 3044 2533 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2493 2956 2533 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2493 2868 2533 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2493 2780 2533 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2493 2692 2533 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2493 2604 2533 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2412 3220 2452 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2412 3132 2452 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2412 3044 2452 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2412 2956 2452 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2412 2868 2452 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2412 2780 2452 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2412 2692 2452 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2412 2604 2452 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2331 3220 2371 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2331 3132 2371 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2331 3044 2371 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2331 2956 2371 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2331 2868 2371 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2331 2780 2371 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2331 2692 2371 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2331 2604 2371 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2250 3220 2290 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2250 3132 2290 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2250 3044 2290 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2250 2956 2290 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2250 2868 2290 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2250 2780 2290 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2250 2692 2290 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2250 2604 2290 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2169 3220 2209 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2169 3132 2209 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2169 3044 2209 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2169 2956 2209 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2169 2868 2209 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2169 2780 2209 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2169 2692 2209 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2169 2604 2209 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2088 3220 2128 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2088 3132 2128 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2088 3044 2128 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2088 2956 2128 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2088 2868 2128 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2088 2780 2128 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2088 2692 2128 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2088 2604 2128 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2007 3220 2047 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2007 3132 2047 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2007 3044 2047 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2007 2956 2047 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2007 2868 2047 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2007 2780 2047 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2007 2692 2047 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 2007 2604 2047 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1926 3220 1966 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1926 3132 1966 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1926 3044 1966 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1926 2956 1966 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1926 2868 1966 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1926 2780 1966 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1926 2692 1966 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1926 2604 1966 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1845 3220 1885 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1845 3132 1885 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1845 3044 1885 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1845 2956 1885 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1845 2868 1885 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1845 2780 1885 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1845 2692 1885 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1845 2604 1885 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1764 3220 1804 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1764 3132 1804 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1764 3044 1804 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1764 2956 1804 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1764 2868 1804 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1764 2780 1804 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1764 2692 1804 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1764 2604 1804 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1683 3220 1723 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1683 3132 1723 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1683 3044 1723 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1683 2956 1723 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1683 2868 1723 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1683 2780 1723 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1683 2692 1723 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1683 2604 1723 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1602 3220 1642 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1602 3132 1642 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1602 3044 1642 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1602 2956 1642 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1602 2868 1642 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1602 2780 1642 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1602 2692 1642 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1602 2604 1642 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1521 3220 1561 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1521 3132 1561 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1521 3044 1561 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1521 2956 1561 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1521 2868 1561 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1521 2780 1561 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1521 2692 1561 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1521 2604 1561 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1440 3220 1480 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1440 3132 1480 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1440 3044 1480 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1440 2956 1480 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1440 2868 1480 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1440 2780 1480 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1440 2692 1480 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1440 2604 1480 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1359 3220 1399 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1359 3132 1399 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1359 3044 1399 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1359 2956 1399 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1359 2868 1399 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1359 2780 1399 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1359 2692 1399 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1359 2604 1399 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1278 3220 1318 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1278 3132 1318 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1278 3044 1318 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1278 2956 1318 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1278 2868 1318 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1278 2780 1318 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1278 2692 1318 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1278 2604 1318 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1197 3220 1237 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1197 3132 1237 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1197 3044 1237 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1197 2956 1237 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1197 2868 1237 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1197 2780 1237 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1197 2692 1237 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1197 2604 1237 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1116 3220 1156 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1116 3132 1156 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1116 3044 1156 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1116 2956 1156 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1116 2868 1156 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1116 2780 1156 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1116 2692 1156 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1116 2604 1156 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1035 3220 1075 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1035 3132 1075 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1035 3044 1075 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1035 2956 1075 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1035 2868 1075 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1035 2780 1075 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1035 2692 1075 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 1035 2604 1075 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 954 3220 994 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 954 3132 994 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 954 3044 994 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 954 2956 994 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 954 2868 994 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 954 2780 994 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 954 2692 994 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 954 2604 994 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 873 3220 913 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 873 3132 913 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 873 3044 913 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 873 2956 913 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 873 2868 913 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 873 2780 913 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 873 2692 913 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 873 2604 913 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 792 3220 832 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 792 3132 832 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 792 3044 832 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 792 2956 832 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 792 2868 832 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 792 2780 832 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 792 2692 832 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 792 2604 832 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 711 3220 751 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 711 3132 751 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 711 3044 751 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 711 2956 751 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 711 2868 751 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 711 2780 751 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 711 2692 751 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 711 2604 751 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 630 3220 670 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 630 3132 670 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 630 3044 670 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 630 2956 670 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 630 2868 670 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 630 2780 670 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 630 2692 670 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 630 2604 670 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 548 3220 588 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 548 3132 588 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 548 3044 588 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 548 2956 588 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 548 2868 588 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 548 2780 588 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 548 2692 588 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 548 2604 588 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 466 3220 506 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 466 3132 506 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 466 3044 506 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 466 2956 506 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 466 2868 506 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 466 2780 506 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 466 2692 506 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 466 2604 506 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 384 3220 424 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 384 3132 424 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 384 3044 424 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 384 2956 424 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 384 2868 424 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 384 2780 424 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 384 2692 424 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 384 2604 424 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 302 3220 342 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 302 3132 342 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 302 3044 342 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 302 2956 342 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 302 2868 342 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 302 2780 342 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 302 2692 342 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 302 2604 342 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 220 3220 260 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 220 3132 260 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 220 3044 260 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 220 2956 260 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 220 2868 260 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 220 2780 260 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 220 2692 260 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 220 2604 260 2644 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 138 3220 178 3260 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 138 3132 178 3172 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 138 3044 178 3084 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 138 2956 178 2996 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 138 2868 178 2908 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 138 2780 178 2820 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 138 2692 178 2732 1 VDDA
port 4 nsew power bidirectional
rlabel via3 s 138 2604 178 2644 1 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 0 13607 254 18600 1 VDDIO
port 6 nsew power bidirectional
rlabel metal4 s 14746 3557 15000 4487 1 VDDIO
port 6 nsew power bidirectional
rlabel metal4 s 14746 13607 15000 18600 1 VDDIO
port 6 nsew power bidirectional
rlabel metal5 s 0 3577 254 4467 1 VDDIO
port 6 nsew power bidirectional
rlabel metal5 s 0 13607 254 18597 1 VDDIO
port 6 nsew power bidirectional
rlabel metal5 s 14746 3577 15000 4467 1 VDDIO
port 6 nsew power bidirectional
rlabel metal5 s 14746 13607 15000 18597 1 VDDIO
port 6 nsew power bidirectional
rlabel metal4 s 14746 12417 15000 13307 1 VDDIO_Q
port 7 nsew power bidirectional
rlabel metal5 s 0 12437 254 13287 1 VDDIO_Q
port 7 nsew power bidirectional
rlabel metal5 s 14746 12437 15000 13287 1 VDDIO_Q
port 7 nsew power bidirectional
rlabel metal4 s 0 9147 254 9213 1 VSSA
port 8 nsew ground bidirectional
rlabel metal4 s 0 9929 254 10165 1 VSSA
port 8 nsew ground bidirectional
rlabel metal4 s 0 10881 254 10947 1 VSSA
port 8 nsew ground bidirectional
rlabel metal4 s 14746 6947 15000 7637 1 VSSA
port 8 nsew ground bidirectional
rlabel metal4 s 14746 9147 15000 9213 1 VSSA
port 8 nsew ground bidirectional
rlabel metal4 s 14746 9929 15000 10165 1 VSSA
port 8 nsew ground bidirectional
rlabel metal4 s 14746 10881 15000 10947 1 VSSA
port 8 nsew ground bidirectional
rlabel metal5 s 0 6968 254 7617 1 VSSA
port 8 nsew ground bidirectional
rlabel metal5 s 0 9147 254 10947 1 VSSA
port 8 nsew ground bidirectional
rlabel metal5 s 14746 6968 15000 7617 1 VSSA
port 8 nsew ground bidirectional
rlabel metal5 s 14746 9147 15000 10947 1 VSSA
port 8 nsew ground bidirectional
rlabel metal4 s 14746 7917 15000 8847 1 VSSD
port 5 nsew ground bidirectional
rlabel metal5 s 0 7937 254 8827 1 VSSD
port 5 nsew ground bidirectional
rlabel metal5 s 14746 7937 15000 8827 1 VSSD
port 5 nsew ground bidirectional
rlabel metal4 s 0 4767 254 5697 1 VSSIO
port 9 nsew ground bidirectional
rlabel metal4 s 14746 34757 15000 39600 1 VSSIO
port 9 nsew ground bidirectional
rlabel metal4 s 14746 4767 15000 5697 1 VSSIO
port 9 nsew ground bidirectional
rlabel metal5 s 0 34757 254 39600 1 VSSIO
port 9 nsew ground bidirectional
rlabel metal5 s 0 4787 254 5677 1 VSSIO
port 9 nsew ground bidirectional
rlabel metal5 s 14746 34757 15000 39600 1 VSSIO
port 9 nsew ground bidirectional
rlabel metal5 s 14746 4787 15000 5677 1 VSSIO
port 9 nsew ground bidirectional
rlabel metal4 s 14746 11247 15000 12137 1 VSSIO_Q
port 10 nsew ground bidirectional
rlabel metal5 s 0 11267 254 12117 1 VSSIO_Q
port 10 nsew ground bidirectional
rlabel metal5 s 14746 11267 15000 12117 1 VSSIO_Q
port 10 nsew ground bidirectional
rlabel metal4 s 14746 5977 15000 6667 1 VSWITCH
port 1 nsew power bidirectional
rlabel metal5 s 0 5997 254 6647 1 VSWITCH
port 1 nsew power bidirectional
rlabel metal5 s 14746 5997 15000 6647 1 VSWITCH
port 1 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 39600
string GDS_END 675976
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 607096
string LEFclass PAD
string LEFsymmetry X Y R90
<< end >>
