magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 1 21 1065 203
rect 30 -17 64 21
<< scnmos >>
rect 81 47 111 177
rect 165 47 195 177
rect 353 47 383 177
rect 437 47 467 177
rect 521 47 551 177
rect 605 47 635 177
rect 705 47 735 177
rect 789 47 819 177
rect 873 47 903 177
rect 957 47 987 177
<< scpmoshvt >>
rect 81 297 111 497
rect 165 297 195 497
rect 353 297 383 497
rect 437 297 467 497
rect 521 297 551 497
rect 605 297 635 497
rect 705 297 735 497
rect 789 297 819 497
rect 873 297 903 497
rect 957 297 987 497
<< ndiff >>
rect 27 163 81 177
rect 27 129 37 163
rect 71 129 81 163
rect 27 95 81 129
rect 27 61 37 95
rect 71 61 81 95
rect 27 47 81 61
rect 111 163 165 177
rect 111 129 121 163
rect 155 129 165 163
rect 111 95 165 129
rect 111 61 121 95
rect 155 61 165 95
rect 111 47 165 61
rect 195 95 353 177
rect 195 61 205 95
rect 239 61 309 95
rect 343 61 353 95
rect 195 47 353 61
rect 383 95 437 177
rect 383 61 393 95
rect 427 61 437 95
rect 383 47 437 61
rect 467 163 521 177
rect 467 129 477 163
rect 511 129 521 163
rect 467 47 521 129
rect 551 95 605 177
rect 551 61 561 95
rect 595 61 605 95
rect 551 47 605 61
rect 635 95 705 177
rect 635 61 654 95
rect 688 61 705 95
rect 635 47 705 61
rect 735 95 789 177
rect 735 61 745 95
rect 779 61 789 95
rect 735 47 789 61
rect 819 163 873 177
rect 819 129 829 163
rect 863 129 873 163
rect 819 47 873 129
rect 903 163 957 177
rect 903 129 913 163
rect 947 129 957 163
rect 903 95 957 129
rect 903 61 913 95
rect 947 61 957 95
rect 903 47 957 61
rect 987 163 1039 177
rect 987 129 997 163
rect 1031 129 1039 163
rect 987 95 1039 129
rect 987 61 997 95
rect 1031 61 1039 95
rect 987 47 1039 61
<< pdiff >>
rect 27 483 81 497
rect 27 449 37 483
rect 71 449 81 483
rect 27 393 81 449
rect 27 359 37 393
rect 71 359 81 393
rect 27 297 81 359
rect 111 409 165 497
rect 111 375 121 409
rect 155 375 165 409
rect 111 341 165 375
rect 111 307 121 341
rect 155 307 165 341
rect 111 297 165 307
rect 195 477 247 497
rect 195 443 205 477
rect 239 443 247 477
rect 195 349 247 443
rect 195 315 205 349
rect 239 315 247 349
rect 195 297 247 315
rect 301 477 353 497
rect 301 443 309 477
rect 343 443 353 477
rect 301 297 353 443
rect 383 409 437 497
rect 383 375 393 409
rect 427 375 437 409
rect 383 297 437 375
rect 467 477 521 497
rect 467 443 477 477
rect 511 443 521 477
rect 467 297 521 443
rect 551 409 605 497
rect 551 375 561 409
rect 595 375 605 409
rect 551 297 605 375
rect 635 477 705 497
rect 635 443 653 477
rect 687 443 705 477
rect 635 407 705 443
rect 635 373 653 407
rect 687 373 705 407
rect 635 297 705 373
rect 735 477 789 497
rect 735 443 745 477
rect 779 443 789 477
rect 735 297 789 443
rect 819 477 873 497
rect 819 443 829 477
rect 863 443 873 477
rect 819 409 873 443
rect 819 375 829 409
rect 863 375 873 409
rect 819 297 873 375
rect 903 477 957 497
rect 903 443 913 477
rect 947 443 957 477
rect 903 297 957 443
rect 987 477 1044 497
rect 987 443 998 477
rect 1032 443 1044 477
rect 987 409 1044 443
rect 987 375 998 409
rect 1032 375 1044 409
rect 987 341 1044 375
rect 987 307 998 341
rect 1032 307 1044 341
rect 987 297 1044 307
<< ndiffc >>
rect 37 129 71 163
rect 37 61 71 95
rect 121 129 155 163
rect 121 61 155 95
rect 205 61 239 95
rect 309 61 343 95
rect 393 61 427 95
rect 477 129 511 163
rect 561 61 595 95
rect 654 61 688 95
rect 745 61 779 95
rect 829 129 863 163
rect 913 129 947 163
rect 913 61 947 95
rect 997 129 1031 163
rect 997 61 1031 95
<< pdiffc >>
rect 37 449 71 483
rect 37 359 71 393
rect 121 375 155 409
rect 121 307 155 341
rect 205 443 239 477
rect 205 315 239 349
rect 309 443 343 477
rect 393 375 427 409
rect 477 443 511 477
rect 561 375 595 409
rect 653 443 687 477
rect 653 373 687 407
rect 745 443 779 477
rect 829 443 863 477
rect 829 375 863 409
rect 913 443 947 477
rect 998 443 1032 477
rect 998 375 1032 409
rect 998 307 1032 341
<< poly >>
rect 81 497 111 523
rect 165 497 195 523
rect 353 497 383 523
rect 437 497 467 523
rect 521 497 551 523
rect 605 497 635 523
rect 705 497 735 523
rect 789 497 819 523
rect 873 497 903 523
rect 957 497 987 523
rect 81 265 111 297
rect 165 265 195 297
rect 353 265 383 297
rect 437 265 467 297
rect 521 265 551 297
rect 605 265 635 297
rect 705 265 735 297
rect 789 265 819 297
rect 873 265 903 297
rect 957 265 987 297
rect 22 249 195 265
rect 22 215 34 249
rect 68 215 195 249
rect 22 199 195 215
rect 341 249 395 265
rect 341 215 351 249
rect 385 215 395 249
rect 341 199 395 215
rect 437 249 551 265
rect 437 215 477 249
rect 511 215 551 249
rect 437 199 551 215
rect 593 249 647 265
rect 593 215 603 249
rect 637 215 647 249
rect 593 199 647 215
rect 693 249 747 265
rect 693 215 703 249
rect 737 215 747 249
rect 693 199 747 215
rect 789 249 903 265
rect 789 215 829 249
rect 863 215 903 249
rect 789 199 903 215
rect 945 249 999 265
rect 945 215 955 249
rect 989 215 999 249
rect 945 199 999 215
rect 81 177 111 199
rect 165 177 195 199
rect 353 177 383 199
rect 437 177 467 199
rect 521 177 551 199
rect 605 177 635 199
rect 705 177 735 199
rect 789 177 819 199
rect 873 177 903 199
rect 957 177 987 199
rect 81 21 111 47
rect 165 21 195 47
rect 353 21 383 47
rect 437 21 467 47
rect 521 21 551 47
rect 605 21 635 47
rect 705 21 735 47
rect 789 21 819 47
rect 873 21 903 47
rect 957 21 987 47
<< polycont >>
rect 34 215 68 249
rect 351 215 385 249
rect 477 215 511 249
rect 603 215 637 249
rect 703 215 737 249
rect 829 215 863 249
rect 955 215 989 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 18 483 255 493
rect 18 449 37 483
rect 71 477 255 483
rect 71 459 205 477
rect 71 449 87 459
rect 18 393 87 449
rect 239 443 255 477
rect 18 359 37 393
rect 71 359 87 393
rect 121 409 171 425
rect 155 375 171 409
rect 121 341 171 375
rect 18 249 84 323
rect 18 215 34 249
rect 68 215 84 249
rect 155 307 171 341
rect 121 181 171 307
rect 205 391 255 443
rect 301 477 695 493
rect 301 443 309 477
rect 343 459 477 477
rect 343 443 351 459
rect 301 425 351 443
rect 469 443 477 459
rect 511 459 653 477
rect 511 443 519 459
rect 469 425 519 443
rect 645 443 653 459
rect 687 443 695 477
rect 385 409 435 425
rect 385 391 393 409
rect 205 375 393 391
rect 427 391 435 409
rect 553 409 603 425
rect 553 391 561 409
rect 427 375 561 391
rect 595 375 603 409
rect 205 357 603 375
rect 645 407 695 443
rect 737 477 787 527
rect 737 443 745 477
rect 779 443 787 477
rect 737 425 787 443
rect 821 477 871 493
rect 821 443 829 477
rect 863 443 871 477
rect 645 373 653 407
rect 687 391 695 407
rect 821 409 871 443
rect 905 477 955 527
rect 905 443 913 477
rect 947 443 955 477
rect 905 425 955 443
rect 998 477 1039 493
rect 1032 443 1039 477
rect 821 391 829 409
rect 687 375 829 391
rect 863 391 871 409
rect 998 409 1039 443
rect 863 375 998 391
rect 1032 375 1039 409
rect 687 373 1039 375
rect 645 357 1039 373
rect 205 349 255 357
rect 239 315 255 349
rect 998 341 1039 357
rect 205 299 255 315
rect 301 289 653 323
rect 301 249 408 289
rect 301 215 351 249
rect 385 215 408 249
rect 442 249 553 255
rect 442 215 477 249
rect 511 215 553 249
rect 587 249 653 289
rect 587 215 603 249
rect 637 215 653 249
rect 687 289 964 323
rect 1032 307 1039 341
rect 998 291 1039 307
rect 687 249 753 289
rect 930 255 964 289
rect 687 215 703 249
rect 737 215 753 249
rect 797 249 896 255
rect 797 215 829 249
rect 863 215 896 249
rect 930 249 1087 255
rect 930 215 955 249
rect 989 215 1087 249
rect 21 163 71 179
rect 121 173 879 181
rect 21 129 37 163
rect 21 95 71 129
rect 21 61 37 95
rect 105 163 879 173
rect 105 129 121 163
rect 155 145 477 163
rect 155 129 171 145
rect 457 129 477 145
rect 511 145 829 163
rect 511 129 527 145
rect 813 129 829 145
rect 863 129 879 163
rect 913 163 963 181
rect 947 129 963 163
rect 105 95 171 129
rect 105 61 121 95
rect 155 61 171 95
rect 205 95 343 111
rect 654 95 688 111
rect 913 95 963 129
rect 239 61 309 95
rect 21 17 71 61
rect 205 17 343 61
rect 377 61 393 95
rect 427 61 561 95
rect 595 61 611 95
rect 377 51 611 61
rect 654 17 688 61
rect 729 61 745 95
rect 779 61 913 95
rect 947 61 963 95
rect 729 51 963 61
rect 997 163 1031 181
rect 997 95 1031 129
rect 997 17 1031 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel locali s 310 289 344 323 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 C1
port 5 nsew signal input
flabel locali s 1046 221 1080 255 0 FreeSans 400 180 0 0 A2
port 2 nsew signal input
flabel locali s 862 221 896 255 0 FreeSans 400 180 0 0 A1
port 1 nsew signal input
flabel locali s 494 221 528 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 310 221 344 255 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 400 0 0 0 Y
port 10 nsew signal output
flabel locali s 30 289 64 323 0 FreeSans 400 0 0 0 C1
port 5 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 a221oi_2
rlabel metal1 s 0 -48 1104 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1104 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_END 3674448
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3665274
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 27.600 0.000 
<< end >>
