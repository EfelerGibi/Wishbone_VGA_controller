magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< pwell >>
rect 251 238 275 289
<< locali >>
rect 0 338 354 354
rect 0 304 16 338
rect 50 304 88 338
rect 122 304 160 338
rect 194 304 232 338
rect 266 304 304 338
rect 338 304 354 338
rect 0 266 354 304
rect 0 232 16 266
rect 50 232 304 266
rect 338 232 354 266
rect 0 194 354 232
rect 0 160 16 194
rect 50 160 304 194
rect 338 160 354 194
rect 0 122 354 160
rect 0 88 16 122
rect 50 88 304 122
rect 338 88 354 122
rect 0 50 354 88
rect 0 16 16 50
rect 50 16 88 50
rect 122 16 160 50
rect 194 16 232 50
rect 266 16 304 50
rect 338 16 354 50
rect 0 0 354 16
<< viali >>
rect 16 304 50 338
rect 88 304 122 338
rect 160 304 194 338
rect 232 304 266 338
rect 304 304 338 338
rect 16 232 50 266
rect 304 232 338 266
rect 16 160 50 194
rect 304 160 338 194
rect 16 88 50 122
rect 304 88 338 122
rect 16 16 50 50
rect 88 16 122 50
rect 160 16 194 50
rect 232 16 266 50
rect 304 16 338 50
<< metal1 >>
rect 0 347 354 354
rect 0 338 64 347
rect 116 338 238 347
rect 290 338 354 347
rect 0 304 16 338
rect 50 304 64 338
rect 122 304 160 338
rect 194 304 232 338
rect 290 304 304 338
rect 338 304 354 338
rect 0 295 64 304
rect 116 295 238 304
rect 290 295 354 304
rect 0 290 354 295
rect 0 238 7 290
rect 59 288 295 290
rect 59 238 66 288
rect 0 232 16 238
rect 50 232 66 238
rect 0 194 66 232
rect 0 160 16 194
rect 50 160 66 194
rect 0 122 66 160
rect 0 116 16 122
rect 50 116 66 122
rect 0 64 7 116
rect 59 66 66 116
rect 94 204 122 260
rect 150 254 204 260
rect 150 204 151 254
rect 94 203 151 204
rect 146 202 151 203
rect 203 204 204 254
rect 232 204 260 260
rect 203 203 260 204
rect 203 202 208 203
rect 146 152 208 202
rect 146 151 151 152
rect 94 150 151 151
rect 94 94 122 150
rect 150 100 151 150
rect 203 151 208 152
rect 203 150 260 151
rect 203 100 204 150
rect 150 94 204 100
rect 232 94 260 150
rect 288 238 295 288
rect 347 238 354 290
rect 288 232 304 238
rect 338 232 354 238
rect 288 194 354 232
rect 288 160 304 194
rect 338 160 354 194
rect 288 122 354 160
rect 288 116 304 122
rect 338 116 354 122
rect 288 66 295 116
rect 59 64 295 66
rect 347 64 354 116
rect 0 59 354 64
rect 0 50 64 59
rect 116 50 238 59
rect 290 50 354 59
rect 0 16 16 50
rect 50 16 64 50
rect 122 16 160 50
rect 194 16 232 50
rect 290 16 304 50
rect 338 16 354 50
rect 0 7 64 16
rect 116 7 238 16
rect 290 7 354 16
rect 0 0 354 7
<< via1 >>
rect 64 338 116 347
rect 238 338 290 347
rect 64 304 88 338
rect 88 304 116 338
rect 238 304 266 338
rect 266 304 290 338
rect 64 295 116 304
rect 238 295 290 304
rect 7 266 59 290
rect 7 238 16 266
rect 16 238 50 266
rect 50 238 59 266
rect 7 88 16 116
rect 16 88 50 116
rect 50 88 59 116
rect 7 64 59 88
rect 94 151 146 203
rect 151 202 203 254
rect 151 100 203 152
rect 208 151 260 203
rect 295 266 347 290
rect 295 238 304 266
rect 304 238 338 266
rect 338 238 347 266
rect 295 88 304 116
rect 304 88 338 116
rect 338 88 347 116
rect 295 64 347 88
rect 64 50 116 59
rect 238 50 290 59
rect 64 16 88 50
rect 88 16 116 50
rect 238 16 266 50
rect 266 16 290 50
rect 64 7 116 16
rect 238 7 290 16
<< metal2 >>
rect 0 347 122 354
rect 0 295 64 347
rect 116 295 122 347
rect 0 290 122 295
rect 0 238 7 290
rect 59 288 122 290
rect 59 238 66 288
rect 150 260 204 354
rect 232 347 354 354
rect 232 295 238 347
rect 290 295 354 347
rect 232 290 354 295
rect 232 288 295 290
rect 0 232 66 238
rect 94 254 260 260
rect 94 232 151 254
rect 150 204 151 232
rect 0 203 151 204
rect 0 151 94 203
rect 146 202 151 203
rect 203 232 260 254
rect 288 238 295 288
rect 347 238 354 290
rect 288 232 354 238
rect 203 204 204 232
rect 203 203 354 204
rect 203 202 208 203
rect 146 152 208 202
rect 146 151 151 152
rect 0 150 151 151
rect 150 122 151 150
rect 0 116 66 122
rect 0 64 7 116
rect 59 66 66 116
rect 94 100 151 122
rect 203 151 208 152
rect 260 151 354 203
rect 203 150 354 151
rect 203 122 204 150
rect 203 100 260 122
rect 94 94 260 100
rect 288 116 354 122
rect 59 64 122 66
rect 0 59 122 64
rect 0 7 64 59
rect 116 7 122 59
rect 0 0 122 7
rect 150 0 204 94
rect 288 66 295 116
rect 232 64 295 66
rect 347 64 354 116
rect 232 59 354 64
rect 232 7 238 59
rect 290 7 354 59
rect 232 0 354 7
<< metal3 >>
rect -211 -211 565 565
<< labels >>
flabel metal3 s 216 157 250 218 0 FreeSans 200 0 0 0 MET3
port 4 nsew
flabel metal2 s 62 307 88 337 0 FreeSans 400 0 0 0 C0
port 1 nsew
flabel metal2 s 160 304 198 341 0 FreeSans 400 0 0 0 C1
port 2 nsew
flabel pwell s 251 238 275 289 0 FreeSans 200 0 0 0 SUB
port 3 nsew
<< properties >>
string GDS_END 59910
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 55686
string device primitive
<< end >>
