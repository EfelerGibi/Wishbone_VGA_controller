magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect 0 0 810 408
<< pmos >>
rect 89 36 119 372
rect 175 36 205 372
rect 261 36 291 372
rect 347 36 377 372
rect 433 36 463 372
rect 519 36 549 372
rect 605 36 635 372
rect 691 36 721 372
<< pdiff >>
rect 36 329 89 372
rect 36 295 44 329
rect 78 295 89 329
rect 36 257 89 295
rect 36 223 44 257
rect 78 223 89 257
rect 36 185 89 223
rect 36 151 44 185
rect 78 151 89 185
rect 36 113 89 151
rect 36 79 44 113
rect 78 79 89 113
rect 36 36 89 79
rect 119 329 175 372
rect 119 295 130 329
rect 164 295 175 329
rect 119 257 175 295
rect 119 223 130 257
rect 164 223 175 257
rect 119 185 175 223
rect 119 151 130 185
rect 164 151 175 185
rect 119 113 175 151
rect 119 79 130 113
rect 164 79 175 113
rect 119 36 175 79
rect 205 329 261 372
rect 205 295 216 329
rect 250 295 261 329
rect 205 257 261 295
rect 205 223 216 257
rect 250 223 261 257
rect 205 185 261 223
rect 205 151 216 185
rect 250 151 261 185
rect 205 113 261 151
rect 205 79 216 113
rect 250 79 261 113
rect 205 36 261 79
rect 291 329 347 372
rect 291 295 302 329
rect 336 295 347 329
rect 291 257 347 295
rect 291 223 302 257
rect 336 223 347 257
rect 291 185 347 223
rect 291 151 302 185
rect 336 151 347 185
rect 291 113 347 151
rect 291 79 302 113
rect 336 79 347 113
rect 291 36 347 79
rect 377 329 433 372
rect 377 295 388 329
rect 422 295 433 329
rect 377 257 433 295
rect 377 223 388 257
rect 422 223 433 257
rect 377 185 433 223
rect 377 151 388 185
rect 422 151 433 185
rect 377 113 433 151
rect 377 79 388 113
rect 422 79 433 113
rect 377 36 433 79
rect 463 329 519 372
rect 463 295 474 329
rect 508 295 519 329
rect 463 257 519 295
rect 463 223 474 257
rect 508 223 519 257
rect 463 185 519 223
rect 463 151 474 185
rect 508 151 519 185
rect 463 113 519 151
rect 463 79 474 113
rect 508 79 519 113
rect 463 36 519 79
rect 549 329 605 372
rect 549 295 560 329
rect 594 295 605 329
rect 549 257 605 295
rect 549 223 560 257
rect 594 223 605 257
rect 549 185 605 223
rect 549 151 560 185
rect 594 151 605 185
rect 549 113 605 151
rect 549 79 560 113
rect 594 79 605 113
rect 549 36 605 79
rect 635 329 691 372
rect 635 295 646 329
rect 680 295 691 329
rect 635 257 691 295
rect 635 223 646 257
rect 680 223 691 257
rect 635 185 691 223
rect 635 151 646 185
rect 680 151 691 185
rect 635 113 691 151
rect 635 79 646 113
rect 680 79 691 113
rect 635 36 691 79
rect 721 329 774 372
rect 721 295 732 329
rect 766 295 774 329
rect 721 257 774 295
rect 721 223 732 257
rect 766 223 774 257
rect 721 185 774 223
rect 721 151 732 185
rect 766 151 774 185
rect 721 113 774 151
rect 721 79 732 113
rect 766 79 774 113
rect 721 36 774 79
<< pdiffc >>
rect 44 295 78 329
rect 44 223 78 257
rect 44 151 78 185
rect 44 79 78 113
rect 130 295 164 329
rect 130 223 164 257
rect 130 151 164 185
rect 130 79 164 113
rect 216 295 250 329
rect 216 223 250 257
rect 216 151 250 185
rect 216 79 250 113
rect 302 295 336 329
rect 302 223 336 257
rect 302 151 336 185
rect 302 79 336 113
rect 388 295 422 329
rect 388 223 422 257
rect 388 151 422 185
rect 388 79 422 113
rect 474 295 508 329
rect 474 223 508 257
rect 474 151 508 185
rect 474 79 508 113
rect 560 295 594 329
rect 560 223 594 257
rect 560 151 594 185
rect 560 79 594 113
rect 646 295 680 329
rect 646 223 680 257
rect 646 151 680 185
rect 646 79 680 113
rect 732 295 766 329
rect 732 223 766 257
rect 732 151 766 185
rect 732 79 766 113
<< poly >>
rect 89 455 721 471
rect 89 421 150 455
rect 184 421 218 455
rect 252 421 286 455
rect 320 421 354 455
rect 388 421 422 455
rect 456 421 490 455
rect 524 421 558 455
rect 592 421 626 455
rect 660 421 721 455
rect 89 398 721 421
rect 89 372 119 398
rect 175 372 205 398
rect 261 372 291 398
rect 347 372 377 398
rect 433 372 463 398
rect 519 372 549 398
rect 605 372 635 398
rect 691 372 721 398
rect 89 10 119 36
rect 175 10 205 36
rect 261 10 291 36
rect 347 10 377 36
rect 433 10 463 36
rect 519 10 549 36
rect 605 10 635 36
rect 691 10 721 36
<< polycont >>
rect 150 421 184 455
rect 218 421 252 455
rect 286 421 320 455
rect 354 421 388 455
rect 422 421 456 455
rect 490 421 524 455
rect 558 421 592 455
rect 626 421 660 455
<< locali >>
rect 134 455 676 471
rect 134 421 136 455
rect 184 421 208 455
rect 252 421 280 455
rect 320 421 352 455
rect 388 421 422 455
rect 458 421 490 455
rect 530 421 558 455
rect 602 421 626 455
rect 674 421 676 455
rect 134 403 676 421
rect 44 329 78 357
rect 44 257 78 295
rect 44 185 78 223
rect 44 113 78 151
rect 44 51 78 79
rect 130 329 164 357
rect 130 257 164 295
rect 130 185 164 223
rect 130 113 164 151
rect 130 51 164 79
rect 216 329 250 357
rect 216 257 250 295
rect 216 185 250 223
rect 216 113 250 151
rect 216 51 250 79
rect 302 329 336 357
rect 302 257 336 295
rect 302 185 336 223
rect 302 113 336 151
rect 302 51 336 79
rect 388 329 422 357
rect 388 257 422 295
rect 388 185 422 223
rect 388 113 422 151
rect 388 51 422 79
rect 474 329 508 357
rect 474 257 508 295
rect 474 185 508 223
rect 474 113 508 151
rect 474 51 508 79
rect 560 329 594 357
rect 560 257 594 295
rect 560 185 594 223
rect 560 113 594 151
rect 560 51 594 79
rect 646 329 680 357
rect 646 257 680 295
rect 646 185 680 223
rect 646 113 680 151
rect 646 51 680 79
rect 732 329 766 357
rect 732 257 766 295
rect 732 185 766 223
rect 732 113 766 151
rect 732 51 766 79
<< viali >>
rect 136 421 150 455
rect 150 421 170 455
rect 208 421 218 455
rect 218 421 242 455
rect 280 421 286 455
rect 286 421 314 455
rect 352 421 354 455
rect 354 421 386 455
rect 424 421 456 455
rect 456 421 458 455
rect 496 421 524 455
rect 524 421 530 455
rect 568 421 592 455
rect 592 421 602 455
rect 640 421 660 455
rect 660 421 674 455
rect 44 295 78 329
rect 44 223 78 257
rect 44 151 78 185
rect 44 79 78 113
rect 130 295 164 329
rect 130 223 164 257
rect 130 151 164 185
rect 130 79 164 113
rect 216 295 250 329
rect 216 223 250 257
rect 216 151 250 185
rect 216 79 250 113
rect 302 295 336 329
rect 302 223 336 257
rect 302 151 336 185
rect 302 79 336 113
rect 388 295 422 329
rect 388 223 422 257
rect 388 151 422 185
rect 388 79 422 113
rect 474 295 508 329
rect 474 223 508 257
rect 474 151 508 185
rect 474 79 508 113
rect 560 295 594 329
rect 560 223 594 257
rect 560 151 594 185
rect 560 79 594 113
rect 646 295 680 329
rect 646 223 680 257
rect 646 151 680 185
rect 646 79 680 113
rect 732 295 766 329
rect 732 223 766 257
rect 732 151 766 185
rect 732 79 766 113
<< metal1 >>
rect 124 455 686 467
rect 124 421 136 455
rect 170 421 208 455
rect 242 421 280 455
rect 314 421 352 455
rect 386 421 424 455
rect 458 421 496 455
rect 530 421 568 455
rect 602 421 640 455
rect 674 421 686 455
rect 124 409 686 421
rect 38 329 84 357
rect 38 295 44 329
rect 78 295 84 329
rect 38 257 84 295
rect 38 223 44 257
rect 78 223 84 257
rect 38 185 84 223
rect 38 151 44 185
rect 78 151 84 185
rect 38 113 84 151
rect 38 79 44 113
rect 78 79 84 113
rect 38 -29 84 79
rect 121 346 173 357
rect 121 282 173 294
rect 121 223 130 230
rect 164 223 173 230
rect 121 185 173 223
rect 121 151 130 185
rect 164 151 173 185
rect 121 113 173 151
rect 121 79 130 113
rect 164 79 173 113
rect 121 51 173 79
rect 210 329 256 357
rect 210 295 216 329
rect 250 295 256 329
rect 210 257 256 295
rect 210 223 216 257
rect 250 223 256 257
rect 210 185 256 223
rect 210 151 216 185
rect 250 151 256 185
rect 210 113 256 151
rect 210 79 216 113
rect 250 79 256 113
rect 210 -29 256 79
rect 293 346 345 357
rect 293 282 345 294
rect 293 223 302 230
rect 336 223 345 230
rect 293 185 345 223
rect 293 151 302 185
rect 336 151 345 185
rect 293 113 345 151
rect 293 79 302 113
rect 336 79 345 113
rect 293 51 345 79
rect 382 329 428 357
rect 382 295 388 329
rect 422 295 428 329
rect 382 257 428 295
rect 382 223 388 257
rect 422 223 428 257
rect 382 185 428 223
rect 382 151 388 185
rect 422 151 428 185
rect 382 113 428 151
rect 382 79 388 113
rect 422 79 428 113
rect 382 -29 428 79
rect 465 346 517 357
rect 465 282 517 294
rect 465 223 474 230
rect 508 223 517 230
rect 465 185 517 223
rect 465 151 474 185
rect 508 151 517 185
rect 465 113 517 151
rect 465 79 474 113
rect 508 79 517 113
rect 465 51 517 79
rect 554 329 600 357
rect 554 295 560 329
rect 594 295 600 329
rect 554 257 600 295
rect 554 223 560 257
rect 594 223 600 257
rect 554 185 600 223
rect 554 151 560 185
rect 594 151 600 185
rect 554 113 600 151
rect 554 79 560 113
rect 594 79 600 113
rect 554 -29 600 79
rect 637 346 689 357
rect 637 282 689 294
rect 637 223 646 230
rect 680 223 689 230
rect 637 185 689 223
rect 637 151 646 185
rect 680 151 689 185
rect 637 113 689 151
rect 637 79 646 113
rect 680 79 689 113
rect 637 51 689 79
rect 726 329 772 357
rect 726 295 732 329
rect 766 295 772 329
rect 726 257 772 295
rect 726 223 732 257
rect 766 223 772 257
rect 726 185 772 223
rect 726 151 732 185
rect 766 151 772 185
rect 726 113 772 151
rect 726 79 732 113
rect 766 79 772 113
rect 726 -29 772 79
rect 38 -89 772 -29
<< via1 >>
rect 121 329 173 346
rect 121 295 130 329
rect 130 295 164 329
rect 164 295 173 329
rect 121 294 173 295
rect 121 257 173 282
rect 121 230 130 257
rect 130 230 164 257
rect 164 230 173 257
rect 293 329 345 346
rect 293 295 302 329
rect 302 295 336 329
rect 336 295 345 329
rect 293 294 345 295
rect 293 257 345 282
rect 293 230 302 257
rect 302 230 336 257
rect 336 230 345 257
rect 465 329 517 346
rect 465 295 474 329
rect 474 295 508 329
rect 508 295 517 329
rect 465 294 517 295
rect 465 257 517 282
rect 465 230 474 257
rect 474 230 508 257
rect 508 230 517 257
rect 637 329 689 346
rect 637 295 646 329
rect 646 295 680 329
rect 680 295 689 329
rect 637 294 689 295
rect 637 257 689 282
rect 637 230 646 257
rect 646 230 680 257
rect 680 230 689 257
<< metal2 >>
rect 114 356 180 365
rect 114 300 119 356
rect 175 300 180 356
rect 114 294 121 300
rect 173 294 180 300
rect 114 282 180 294
rect 114 276 121 282
rect 173 276 180 282
rect 114 220 119 276
rect 175 220 180 276
rect 114 211 180 220
rect 286 356 352 365
rect 286 300 291 356
rect 347 300 352 356
rect 286 294 293 300
rect 345 294 352 300
rect 286 282 352 294
rect 286 276 293 282
rect 345 276 352 282
rect 286 220 291 276
rect 347 220 352 276
rect 286 211 352 220
rect 458 356 524 365
rect 458 300 463 356
rect 519 300 524 356
rect 458 294 465 300
rect 517 294 524 300
rect 458 282 524 294
rect 458 276 465 282
rect 517 276 524 282
rect 458 220 463 276
rect 519 220 524 276
rect 458 211 524 220
rect 630 356 696 365
rect 630 300 635 356
rect 691 300 696 356
rect 630 294 637 300
rect 689 294 696 300
rect 630 282 696 294
rect 630 276 637 282
rect 689 276 696 282
rect 630 220 635 276
rect 691 220 696 276
rect 630 211 696 220
<< via2 >>
rect 119 346 175 356
rect 119 300 121 346
rect 121 300 173 346
rect 173 300 175 346
rect 119 230 121 276
rect 121 230 173 276
rect 173 230 175 276
rect 119 220 175 230
rect 291 346 347 356
rect 291 300 293 346
rect 293 300 345 346
rect 345 300 347 346
rect 291 230 293 276
rect 293 230 345 276
rect 345 230 347 276
rect 291 220 347 230
rect 463 346 519 356
rect 463 300 465 346
rect 465 300 517 346
rect 517 300 519 346
rect 463 230 465 276
rect 465 230 517 276
rect 517 230 519 276
rect 463 220 519 230
rect 635 346 691 356
rect 635 300 637 346
rect 637 300 689 346
rect 689 300 691 346
rect 635 230 637 276
rect 637 230 689 276
rect 689 230 691 276
rect 635 220 691 230
<< metal3 >>
rect 114 356 696 365
rect 114 300 119 356
rect 175 300 291 356
rect 347 300 463 356
rect 519 300 635 356
rect 691 300 696 356
rect 114 299 696 300
rect 114 276 180 299
rect 114 220 119 276
rect 175 220 180 276
rect 114 211 180 220
rect 286 276 352 299
rect 286 220 291 276
rect 347 220 352 276
rect 286 211 352 220
rect 458 276 524 299
rect 458 220 463 276
rect 519 220 524 276
rect 458 211 524 220
rect 630 276 696 299
rect 630 220 635 276
rect 691 220 696 276
rect 630 211 696 220
<< labels >>
flabel metal3 s 114 299 696 365 0 FreeSans 400 0 0 0 DRAIN
port 2 nsew
flabel metal1 s 124 409 686 467 0 FreeSans 400 0 0 0 GATE
port 3 nsew
flabel metal1 s 38 -89 772 -29 0 FreeSans 400 0 0 0 SOURCE
port 4 nsew
flabel nwell s 83 400 86 405 0 FreeSans 400 0 0 0 BULK
port 5 nsew
<< properties >>
string GDS_END 9275288
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9261312
string path 1.525 8.925 1.525 -2.225 
<< end >>
