magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1 201 1637 203
rect 1 23 1951 201
rect 1 21 479 23
rect 956 21 1140 23
rect 1552 21 1951 23
rect 47 -17 81 21
<< locali >>
rect 139 409 173 493
rect 307 409 341 493
rect 139 291 341 409
rect 139 288 284 291
rect 221 185 284 288
rect 119 166 307 185
rect 119 132 321 166
rect 119 70 153 132
rect 287 70 321 132
rect 576 199 703 265
rect 1541 289 1657 323
rect 1541 199 1575 289
rect 1705 215 1787 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 55 427 89 527
rect 207 443 273 527
rect 375 443 441 527
rect 475 447 783 481
rect 826 447 907 481
rect 941 447 1007 527
rect 1074 455 1693 489
rect 1783 455 1849 527
rect 475 409 509 447
rect 873 413 907 447
rect 1074 413 1108 455
rect 375 375 509 409
rect 578 379 839 413
rect 873 379 1108 413
rect 375 265 409 375
rect 474 307 771 341
rect 364 193 409 265
rect 375 173 409 193
rect 375 139 473 173
rect 35 17 69 109
rect 187 17 253 93
rect 371 17 405 105
rect 439 85 473 139
rect 508 119 542 307
rect 737 265 771 307
rect 805 339 839 379
rect 805 305 911 339
rect 854 275 911 305
rect 737 199 811 265
rect 598 131 820 165
rect 682 85 752 91
rect 439 51 752 85
rect 786 85 820 131
rect 854 119 888 275
rect 945 241 979 379
rect 1025 289 1108 343
rect 922 210 979 241
rect 922 209 978 210
rect 922 208 976 209
rect 922 207 973 208
rect 922 85 956 207
rect 786 51 956 85
rect 990 17 1024 177
rect 1060 83 1108 289
rect 1143 119 1177 421
rect 1215 178 1249 455
rect 1883 421 1935 493
rect 1283 323 1366 409
rect 1473 387 1935 421
rect 1283 289 1439 323
rect 1286 199 1371 254
rect 1215 165 1255 178
rect 1215 144 1294 165
rect 1221 131 1294 144
rect 1143 97 1187 119
rect 1143 53 1226 97
rect 1260 64 1294 131
rect 1328 126 1371 199
rect 1405 85 1439 289
rect 1473 119 1507 387
rect 1838 375 1935 387
rect 1691 299 1855 341
rect 1821 265 1855 299
rect 1609 189 1671 255
rect 1821 199 1867 265
rect 1609 146 1650 189
rect 1821 181 1855 199
rect 1707 150 1855 181
rect 1699 147 1855 150
rect 1541 85 1634 93
rect 1405 51 1634 85
rect 1699 59 1757 147
rect 1901 117 1935 375
rect 1799 17 1833 113
rect 1883 51 1935 117
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< obsm1 >>
rect 865 320 923 329
rect 1325 320 1383 329
rect 865 292 1383 320
rect 865 283 923 292
rect 1325 283 1383 292
rect 1049 184 1107 193
rect 1325 184 1383 193
rect 1601 184 1659 193
rect 1049 156 1659 184
rect 1049 147 1107 156
rect 1325 147 1383 156
rect 1601 147 1659 156
rect 1141 116 1199 125
rect 1693 116 1751 125
rect 1141 88 1751 116
rect 1141 79 1199 88
rect 1693 79 1751 88
<< labels >>
rlabel locali s 1705 215 1787 265 6 A
port 1 nsew signal input
rlabel locali s 1541 199 1575 289 6 B
port 2 nsew signal input
rlabel locali s 1541 289 1657 323 6 B
port 2 nsew signal input
rlabel locali s 576 199 703 265 6 C
port 3 nsew signal input
rlabel metal1 s 0 -48 2024 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 47 -17 81 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1552 21 1951 23 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 956 21 1140 23 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 479 23 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 23 1951 201 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 201 1637 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 2062 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 2024 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 287 70 321 132 6 X
port 8 nsew signal output
rlabel locali s 119 70 153 132 6 X
port 8 nsew signal output
rlabel locali s 119 132 321 166 6 X
port 8 nsew signal output
rlabel locali s 119 166 307 185 6 X
port 8 nsew signal output
rlabel locali s 221 185 284 288 6 X
port 8 nsew signal output
rlabel locali s 139 288 284 291 6 X
port 8 nsew signal output
rlabel locali s 139 291 341 409 6 X
port 8 nsew signal output
rlabel locali s 307 409 341 493 6 X
port 8 nsew signal output
rlabel locali s 139 409 173 493 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2024 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 698948
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 685650
<< end >>
