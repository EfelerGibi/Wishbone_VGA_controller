magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< locali >>
rect 181 742 193 776
rect 227 742 265 776
rect 299 742 337 776
rect 371 742 383 776
rect 181 30 193 64
rect 227 30 265 64
rect 299 30 337 64
rect 371 30 383 64
<< viali >>
rect 193 742 227 776
rect 265 742 299 776
rect 337 742 371 776
rect 193 30 227 64
rect 265 30 299 64
rect 337 30 371 64
<< obsli1 >>
rect 48 672 82 674
rect 48 600 82 638
rect 48 528 82 566
rect 48 456 82 494
rect 48 384 82 422
rect 48 312 82 350
rect 48 240 82 278
rect 48 168 82 206
rect 48 132 82 134
rect 159 98 193 708
rect 265 98 299 708
rect 371 98 405 708
rect 482 672 516 674
rect 482 600 516 638
rect 482 528 516 566
rect 482 456 516 494
rect 482 384 516 422
rect 482 312 516 350
rect 482 240 516 278
rect 482 168 516 206
rect 482 132 516 134
<< obsli1c >>
rect 48 638 82 672
rect 48 566 82 600
rect 48 494 82 528
rect 48 422 82 456
rect 48 350 82 384
rect 48 278 82 312
rect 48 206 82 240
rect 48 134 82 168
rect 482 638 516 672
rect 482 566 516 600
rect 482 494 516 528
rect 482 422 516 456
rect 482 350 516 384
rect 482 278 516 312
rect 482 206 516 240
rect 482 134 516 168
<< metal1 >>
rect 181 776 383 796
rect 181 742 193 776
rect 227 742 265 776
rect 299 742 337 776
rect 371 742 383 776
rect 181 730 383 742
rect 36 672 94 684
rect 36 638 48 672
rect 82 638 94 672
rect 36 600 94 638
rect 36 566 48 600
rect 82 566 94 600
rect 36 528 94 566
rect 36 494 48 528
rect 82 494 94 528
rect 36 456 94 494
rect 36 422 48 456
rect 82 422 94 456
rect 36 384 94 422
rect 36 350 48 384
rect 82 350 94 384
rect 36 312 94 350
rect 36 278 48 312
rect 82 278 94 312
rect 36 240 94 278
rect 36 206 48 240
rect 82 206 94 240
rect 36 168 94 206
rect 36 134 48 168
rect 82 134 94 168
rect 36 122 94 134
rect 470 672 528 684
rect 470 638 482 672
rect 516 638 528 672
rect 470 600 528 638
rect 470 566 482 600
rect 516 566 528 600
rect 470 528 528 566
rect 470 494 482 528
rect 516 494 528 528
rect 470 456 528 494
rect 470 422 482 456
rect 516 422 528 456
rect 470 384 528 422
rect 470 350 482 384
rect 516 350 528 384
rect 470 312 528 350
rect 470 278 482 312
rect 516 278 528 312
rect 470 240 528 278
rect 470 206 482 240
rect 516 206 528 240
rect 470 168 528 206
rect 470 134 482 168
rect 516 134 528 168
rect 470 122 528 134
rect 181 64 383 76
rect 181 30 193 64
rect 227 30 265 64
rect 299 30 337 64
rect 371 30 383 64
rect 181 10 383 30
<< obsm1 >>
rect 150 122 202 684
rect 256 122 308 684
rect 362 122 414 684
<< metal2 >>
rect 10 428 554 684
rect 10 122 554 378
<< labels >>
rlabel metal2 s 10 428 554 684 6 DRAIN
port 1 nsew
rlabel viali s 337 742 371 776 6 GATE
port 2 nsew
rlabel viali s 337 30 371 64 6 GATE
port 2 nsew
rlabel viali s 265 742 299 776 6 GATE
port 2 nsew
rlabel viali s 265 30 299 64 6 GATE
port 2 nsew
rlabel viali s 193 742 227 776 6 GATE
port 2 nsew
rlabel viali s 193 30 227 64 6 GATE
port 2 nsew
rlabel locali s 181 742 383 776 6 GATE
port 2 nsew
rlabel locali s 181 30 383 64 6 GATE
port 2 nsew
rlabel metal1 s 181 730 383 796 6 GATE
port 2 nsew
rlabel metal1 s 181 10 383 76 6 GATE
port 2 nsew
rlabel metal2 s 10 122 554 378 6 SOURCE
port 3 nsew
rlabel metal1 s 36 122 94 684 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 470 122 528 684 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 10 10 554 796
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4949032
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 4938168
<< end >>
