magic
tech sky130A
magscale 1 2
timestamp 1683767628
use sky130_fd_pr__nfet_01v8__example_55959141808575  sky130_fd_pr__nfet_01v8__example_55959141808575_0
timestamp 1683767628
transform 1 0 119 0 1 36
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808574  sky130_fd_pr__pfet_01v8__example_55959141808574_0
timestamp 1683767628
transform 1 0 119 0 -1 682
box -1 0 101 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1683767628
transform -1 0 205 0 -1 349
box 0 0 1 1
<< properties >>
string GDS_END 8126600
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8126166
<< end >>
