magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 273 157 457 201
rect 1673 181 1857 203
rect 1390 157 1857 181
rect 1 21 1857 157
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 175
rect 446 47 476 119
rect 556 47 586 119
rect 652 47 682 131
rect 766 47 796 131
rect 838 47 868 131
rect 1026 47 1056 131
rect 1098 47 1128 131
rect 1194 47 1224 131
rect 1266 47 1296 131
rect 1342 47 1372 131
rect 1466 47 1496 155
rect 1654 47 1684 131
rect 1749 47 1779 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 329 381 497
rect 448 413 478 497
rect 532 413 562 497
rect 652 413 682 497
rect 758 413 788 497
rect 842 413 872 497
rect 926 413 956 497
rect 1002 413 1032 497
rect 1110 413 1140 497
rect 1182 413 1212 497
rect 1370 413 1400 497
rect 1466 329 1496 497
rect 1654 369 1684 497
rect 1749 297 1779 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 93 351 175
rect 299 59 307 93
rect 341 59 351 93
rect 299 47 351 59
rect 381 119 431 175
rect 1416 131 1466 155
rect 601 119 652 131
rect 381 111 446 119
rect 381 77 391 111
rect 425 77 446 111
rect 381 47 446 77
rect 476 93 556 119
rect 476 59 501 93
rect 535 59 556 93
rect 476 47 556 59
rect 586 47 652 119
rect 682 89 766 131
rect 682 55 722 89
rect 756 55 766 89
rect 682 47 766 55
rect 796 47 838 131
rect 868 109 920 131
rect 868 75 878 109
rect 912 75 920 109
rect 868 47 920 75
rect 974 93 1026 131
rect 974 59 982 93
rect 1016 59 1026 93
rect 974 47 1026 59
rect 1056 47 1098 131
rect 1128 95 1194 131
rect 1128 61 1144 95
rect 1178 61 1194 95
rect 1128 47 1194 61
rect 1224 47 1266 131
rect 1296 47 1342 131
rect 1372 113 1466 131
rect 1372 79 1402 113
rect 1436 79 1466 113
rect 1372 47 1466 79
rect 1496 120 1548 155
rect 1699 131 1749 177
rect 1496 86 1506 120
rect 1540 86 1548 120
rect 1496 47 1548 86
rect 1602 119 1654 131
rect 1602 85 1610 119
rect 1644 85 1654 119
rect 1602 47 1654 85
rect 1684 93 1749 131
rect 1684 59 1705 93
rect 1739 59 1749 93
rect 1684 47 1749 59
rect 1779 143 1831 177
rect 1779 109 1789 143
rect 1823 109 1831 143
rect 1779 47 1831 109
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 461 351 497
rect 299 427 307 461
rect 341 427 351 461
rect 299 329 351 427
rect 381 477 448 497
rect 381 443 391 477
rect 425 443 448 477
rect 381 413 448 443
rect 478 484 532 497
rect 478 450 488 484
rect 522 450 532 484
rect 478 413 532 450
rect 562 413 652 497
rect 682 485 758 497
rect 682 451 702 485
rect 736 451 758 485
rect 682 413 758 451
rect 788 459 842 497
rect 788 425 798 459
rect 832 425 842 459
rect 788 413 842 425
rect 872 485 926 497
rect 872 451 882 485
rect 916 451 926 485
rect 872 413 926 451
rect 956 413 1002 497
rect 1032 483 1110 497
rect 1032 449 1042 483
rect 1076 449 1110 483
rect 1032 413 1110 449
rect 1140 413 1182 497
rect 1212 485 1264 497
rect 1212 451 1222 485
rect 1256 451 1264 485
rect 1212 413 1264 451
rect 1318 459 1370 497
rect 1318 425 1326 459
rect 1360 425 1370 459
rect 1318 413 1370 425
rect 1400 459 1466 497
rect 1400 425 1422 459
rect 1456 425 1466 459
rect 1400 413 1466 425
rect 381 409 433 413
rect 381 375 391 409
rect 425 375 433 409
rect 381 329 433 375
rect 1415 329 1466 413
rect 1496 459 1548 497
rect 1496 425 1506 459
rect 1540 425 1548 459
rect 1496 391 1548 425
rect 1496 357 1506 391
rect 1540 357 1548 391
rect 1602 485 1654 497
rect 1602 451 1610 485
rect 1644 451 1654 485
rect 1602 417 1654 451
rect 1602 383 1610 417
rect 1644 383 1654 417
rect 1602 369 1654 383
rect 1684 485 1749 497
rect 1684 451 1705 485
rect 1739 451 1749 485
rect 1684 417 1749 451
rect 1684 383 1705 417
rect 1739 383 1749 417
rect 1684 369 1749 383
rect 1496 329 1548 357
rect 1699 297 1749 369
rect 1779 449 1831 497
rect 1779 415 1789 449
rect 1823 415 1831 449
rect 1779 381 1831 415
rect 1779 347 1789 381
rect 1823 347 1831 381
rect 1779 297 1831 347
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 59 341 93
rect 391 77 425 111
rect 501 59 535 93
rect 722 55 756 89
rect 878 75 912 109
rect 982 59 1016 93
rect 1144 61 1178 95
rect 1402 79 1436 113
rect 1506 86 1540 120
rect 1610 85 1644 119
rect 1705 59 1739 93
rect 1789 109 1823 143
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 427 341 461
rect 391 443 425 477
rect 488 450 522 484
rect 702 451 736 485
rect 798 425 832 459
rect 882 451 916 485
rect 1042 449 1076 483
rect 1222 451 1256 485
rect 1326 425 1360 459
rect 1422 425 1456 459
rect 391 375 425 409
rect 1506 425 1540 459
rect 1506 357 1540 391
rect 1610 451 1644 485
rect 1610 383 1644 417
rect 1705 451 1739 485
rect 1705 383 1739 417
rect 1789 415 1823 449
rect 1789 347 1823 381
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 448 497 478 523
rect 532 497 562 523
rect 652 497 682 523
rect 758 497 788 523
rect 842 497 872 523
rect 926 497 956 523
rect 1002 497 1032 523
rect 1110 497 1140 523
rect 1182 497 1212 523
rect 1370 497 1400 523
rect 1466 497 1496 523
rect 1654 497 1684 523
rect 1749 497 1779 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 280 76 318
rect 22 264 76 280
rect 163 274 193 363
rect 22 230 32 264
rect 66 230 76 264
rect 22 214 76 230
rect 118 264 193 274
rect 351 267 381 329
rect 448 279 478 413
rect 532 375 562 413
rect 652 381 682 413
rect 520 365 586 375
rect 520 331 536 365
rect 570 331 586 365
rect 520 321 586 331
rect 652 365 716 381
rect 652 331 672 365
rect 706 331 716 365
rect 652 315 716 331
rect 118 230 134 264
rect 168 230 193 264
rect 118 220 193 230
rect 46 176 76 214
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 344 251 398 267
rect 344 217 354 251
rect 388 217 398 251
rect 448 249 586 279
rect 344 201 398 217
rect 556 219 586 249
rect 351 175 381 201
rect 446 191 514 207
rect 446 157 470 191
rect 504 157 514 191
rect 446 141 514 157
rect 556 203 610 219
rect 556 169 566 203
rect 600 169 610 203
rect 556 153 610 169
rect 446 119 476 141
rect 556 119 586 153
rect 652 131 682 315
rect 758 229 788 413
rect 842 313 872 413
rect 926 313 956 413
rect 1002 375 1032 413
rect 1002 365 1068 375
rect 1002 331 1018 365
rect 1052 331 1068 365
rect 1002 321 1068 331
rect 830 297 956 313
rect 830 263 840 297
rect 874 263 956 297
rect 1110 291 1140 413
rect 1098 279 1140 291
rect 830 247 956 263
rect 1034 269 1140 279
rect 728 213 788 229
rect 728 179 738 213
rect 772 193 788 213
rect 772 179 796 193
rect 728 163 796 179
rect 766 131 796 163
rect 838 183 868 247
rect 1034 235 1050 269
rect 1084 261 1140 269
rect 1182 365 1212 413
rect 1182 349 1246 365
rect 1182 315 1202 349
rect 1236 315 1246 349
rect 1370 337 1400 413
rect 1182 291 1246 315
rect 1366 307 1400 337
rect 1182 261 1296 291
rect 1084 235 1128 261
rect 1034 225 1128 235
rect 838 147 1056 183
rect 838 131 868 147
rect 1026 131 1056 147
rect 1098 131 1128 225
rect 1170 203 1224 219
rect 1170 169 1180 203
rect 1214 169 1224 203
rect 1170 153 1224 169
rect 1194 131 1224 153
rect 1266 131 1296 261
rect 1366 229 1396 307
rect 1466 285 1496 329
rect 1654 285 1684 369
rect 1342 213 1396 229
rect 1438 269 1684 285
rect 1438 235 1448 269
rect 1482 235 1684 269
rect 1749 265 1779 297
rect 1438 219 1684 235
rect 1342 179 1352 213
rect 1386 179 1396 213
rect 1342 163 1396 179
rect 1342 131 1372 163
rect 1466 155 1496 219
rect 1654 131 1684 219
rect 1726 249 1780 265
rect 1726 215 1736 249
rect 1770 215 1780 249
rect 1726 199 1780 215
rect 1749 177 1779 199
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 446 21 476 47
rect 556 21 586 47
rect 652 21 682 47
rect 766 21 796 47
rect 838 21 868 47
rect 1026 21 1056 47
rect 1098 21 1128 47
rect 1194 21 1224 47
rect 1266 21 1296 47
rect 1342 21 1372 47
rect 1466 21 1496 47
rect 1654 21 1684 47
rect 1749 21 1779 47
<< polycont >>
rect 32 230 66 264
rect 536 331 570 365
rect 672 331 706 365
rect 134 230 168 264
rect 354 217 388 251
rect 470 157 504 191
rect 566 169 600 203
rect 1018 331 1052 365
rect 840 263 874 297
rect 738 179 772 213
rect 1050 235 1084 269
rect 1202 315 1236 349
rect 1180 169 1214 203
rect 1448 235 1482 269
rect 1352 179 1386 213
rect 1736 215 1770 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 237 443 248 477
rect 203 409 248 443
rect 291 461 357 527
rect 291 427 307 461
rect 341 427 357 461
rect 391 477 425 493
rect 686 485 762 527
rect 472 450 488 484
rect 522 450 638 484
rect 686 451 702 485
rect 736 451 762 485
rect 866 485 932 527
rect 798 459 832 475
rect 69 391 168 393
rect 69 375 122 391
rect 35 359 122 375
rect 156 357 168 391
rect 18 264 88 325
rect 18 230 32 264
rect 66 230 88 264
rect 18 195 88 230
rect 122 264 168 357
rect 122 230 134 264
rect 122 161 168 230
rect 35 127 168 161
rect 237 375 248 409
rect 391 409 425 443
rect 203 187 248 375
rect 203 153 214 187
rect 35 119 69 127
rect 203 119 248 153
rect 286 375 391 393
rect 286 359 425 375
rect 286 165 320 359
rect 470 357 494 391
rect 528 365 570 391
rect 528 357 536 365
rect 470 331 536 357
rect 354 251 436 325
rect 388 217 436 251
rect 354 201 436 217
rect 470 315 570 331
rect 470 191 514 315
rect 604 281 638 450
rect 866 451 882 485
rect 916 451 932 485
rect 1188 485 1272 527
rect 1026 449 1042 483
rect 1076 449 1152 483
rect 1188 451 1222 485
rect 1256 451 1272 485
rect 1312 459 1360 475
rect 1026 433 1152 449
rect 798 417 832 425
rect 1118 417 1152 433
rect 1312 425 1326 459
rect 1312 417 1360 425
rect 672 367 946 417
rect 672 365 722 367
rect 706 331 722 365
rect 672 315 722 331
rect 824 297 874 313
rect 824 281 840 297
rect 604 263 840 281
rect 604 247 874 263
rect 604 239 688 247
rect 286 127 425 165
rect 504 157 514 191
rect 470 141 514 157
rect 550 169 566 203
rect 600 187 620 203
rect 550 153 586 169
rect 550 129 620 153
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 237 85 248 119
rect 391 111 425 127
rect 203 69 248 85
rect 103 17 169 59
rect 291 59 307 93
rect 341 59 357 93
rect 654 93 688 239
rect 908 213 946 367
rect 722 179 738 213
rect 772 187 804 213
rect 722 153 770 179
rect 722 147 804 153
rect 862 145 946 213
rect 980 391 1084 393
rect 980 365 1050 391
rect 980 331 1018 365
rect 1052 331 1084 357
rect 1118 383 1360 417
rect 1406 459 1472 527
rect 1696 485 1753 527
rect 1406 425 1422 459
rect 1456 425 1472 459
rect 1406 389 1472 425
rect 1506 459 1540 475
rect 1506 391 1540 425
rect 980 179 1014 331
rect 1048 269 1084 295
rect 1048 221 1050 269
rect 1118 281 1152 383
rect 1594 451 1610 485
rect 1644 451 1660 485
rect 1594 417 1660 451
rect 1594 383 1610 417
rect 1644 383 1660 417
rect 1506 353 1540 357
rect 1506 349 1570 353
rect 1186 315 1202 349
rect 1236 315 1570 349
rect 1118 269 1498 281
rect 1118 247 1448 269
rect 1048 213 1084 221
rect 1164 179 1180 203
rect 980 169 1180 179
rect 1214 169 1230 203
rect 980 145 1230 169
rect 862 109 912 145
rect 391 61 425 77
rect 291 17 357 59
rect 485 59 501 93
rect 535 59 688 93
rect 485 53 688 59
rect 722 89 804 105
rect 756 55 804 89
rect 862 75 878 109
rect 862 59 912 75
rect 952 93 1016 109
rect 1264 95 1298 247
rect 1432 235 1448 247
rect 1482 235 1498 269
rect 1336 179 1352 213
rect 1386 201 1402 213
rect 1386 187 1468 201
rect 1386 179 1422 187
rect 1336 153 1422 179
rect 1456 153 1468 187
rect 1336 147 1468 153
rect 1532 136 1570 315
rect 1506 120 1570 136
rect 952 59 982 93
rect 1128 61 1144 95
rect 1178 61 1298 95
rect 1338 79 1402 113
rect 1436 79 1470 113
rect 722 17 804 55
rect 952 17 1016 59
rect 1338 17 1470 79
rect 1540 86 1570 120
rect 1506 70 1570 86
rect 1610 265 1660 383
rect 1696 451 1705 485
rect 1739 451 1753 485
rect 1696 417 1753 451
rect 1696 383 1705 417
rect 1739 383 1753 417
rect 1696 367 1753 383
rect 1789 449 1840 465
rect 1823 415 1840 449
rect 1789 381 1840 415
rect 1823 347 1840 381
rect 1789 331 1840 347
rect 1610 249 1770 265
rect 1610 215 1736 249
rect 1610 199 1770 215
rect 1610 119 1660 199
rect 1804 159 1840 331
rect 1644 85 1660 119
rect 1789 143 1840 159
rect 1823 109 1840 143
rect 1610 69 1660 85
rect 1696 93 1753 109
rect 1696 59 1705 93
rect 1739 59 1753 93
rect 1696 17 1753 59
rect 1789 53 1840 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 122 357 156 391
rect 214 153 248 187
rect 494 357 528 391
rect 586 169 600 187
rect 600 169 620 187
rect 586 153 620 169
rect 770 179 772 187
rect 772 179 804 187
rect 770 153 804 179
rect 1050 365 1084 391
rect 1050 357 1052 365
rect 1052 357 1084 365
rect 1050 235 1084 255
rect 1050 221 1084 235
rect 1422 153 1456 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 110 391 168 397
rect 110 357 122 391
rect 156 388 168 391
rect 482 391 540 397
rect 482 388 494 391
rect 156 360 494 388
rect 156 357 168 360
rect 110 351 168 357
rect 482 357 494 360
rect 528 388 540 391
rect 1038 391 1096 397
rect 1038 388 1050 391
rect 528 360 1050 388
rect 528 357 540 360
rect 482 351 540 357
rect 1038 357 1050 360
rect 1084 357 1096 391
rect 1038 351 1096 357
rect 1038 255 1096 261
rect 1038 252 1050 255
rect 589 224 1050 252
rect 589 193 632 224
rect 1038 221 1050 224
rect 1084 221 1096 255
rect 1038 215 1096 221
rect 202 187 260 193
rect 202 153 214 187
rect 248 184 260 187
rect 574 187 632 193
rect 574 184 586 187
rect 248 156 586 184
rect 248 153 260 156
rect 202 147 260 153
rect 574 153 586 156
rect 620 153 632 187
rect 574 147 632 153
rect 758 187 816 193
rect 758 153 770 187
rect 804 184 816 187
rect 1410 187 1468 193
rect 1410 184 1422 187
rect 804 156 1422 184
rect 804 153 816 156
rect 758 147 816 153
rect 1410 153 1422 156
rect 1456 153 1468 187
rect 1410 147 1468 153
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
flabel locali s 402 289 436 323 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 402 221 436 255 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 29 527 63 561 3 FreeSans 400 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 1794 425 1828 459 0 FreeSans 400 0 0 0 Q
port 8 nsew signal output
flabel locali s 1794 357 1828 391 0 FreeSans 400 0 0 0 Q
port 8 nsew signal output
flabel locali s 1794 85 1828 119 0 FreeSans 400 0 0 0 Q
port 8 nsew signal output
flabel locali s 770 153 804 187 0 FreeSans 400 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 30 289 64 323 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 29 -17 63 17 3 FreeSans 400 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel nwell s 46 544 46 544 3 FreeSans 400 0 0 0 VPB
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel pwell s 46 0 46 0 3 FreeSans 400 0 0 0 VNB
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 dfstp_1
rlabel locali s 1336 201 1402 213 1 SET_B
port 3 nsew signal input
rlabel locali s 1336 147 1468 201 1 SET_B
port 3 nsew signal input
rlabel metal1 s 1410 184 1468 193 1 SET_B
port 3 nsew signal input
rlabel metal1 s 1410 147 1468 156 1 SET_B
port 3 nsew signal input
rlabel metal1 s 758 184 816 193 1 SET_B
port 3 nsew signal input
rlabel metal1 s 758 156 1468 184 1 SET_B
port 3 nsew signal input
rlabel metal1 s 758 147 816 156 1 SET_B
port 3 nsew signal input
rlabel metal1 s 0 -48 1932 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1932 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1932 544
string GDS_END 2546124
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2530582
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
