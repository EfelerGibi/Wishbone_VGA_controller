magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 833 157 1287 203
rect 1 21 1287 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 435 47 465 131
rect 530 47 560 119
rect 628 47 658 119
rect 723 47 753 131
rect 911 47 941 177
rect 995 47 1025 177
rect 1095 47 1125 177
rect 1179 47 1209 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 369 381 497
rect 435 369 465 497
rect 531 413 561 497
rect 615 413 645 497
rect 711 413 741 497
rect 908 297 938 497
rect 992 297 1022 497
rect 1088 297 1118 497
rect 1179 297 1209 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 119 351 131
rect 299 85 307 119
rect 341 85 351 119
rect 299 47 351 85
rect 381 89 435 131
rect 381 55 391 89
rect 425 55 435 89
rect 381 47 435 55
rect 465 119 515 131
rect 859 165 911 177
rect 859 131 867 165
rect 901 131 911 165
rect 673 119 723 131
rect 465 47 530 119
rect 560 107 628 119
rect 560 73 579 107
rect 613 73 628 107
rect 560 47 628 73
rect 658 47 723 119
rect 753 106 805 131
rect 753 72 763 106
rect 797 72 805 106
rect 753 47 805 72
rect 859 97 911 131
rect 859 63 867 97
rect 901 63 911 97
rect 859 47 911 63
rect 941 47 995 177
rect 1025 89 1095 177
rect 1025 55 1035 89
rect 1069 55 1095 89
rect 1025 47 1095 55
rect 1125 89 1179 177
rect 1125 55 1135 89
rect 1169 55 1179 89
rect 1125 47 1179 55
rect 1209 93 1261 177
rect 1209 59 1219 93
rect 1253 59 1261 93
rect 1209 47 1261 59
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 483 351 497
rect 299 449 307 483
rect 341 449 351 483
rect 299 415 351 449
rect 299 381 307 415
rect 341 381 351 415
rect 299 369 351 381
rect 381 485 435 497
rect 381 451 391 485
rect 425 451 435 485
rect 381 417 435 451
rect 381 383 391 417
rect 425 383 435 417
rect 381 369 435 383
rect 465 413 531 497
rect 561 485 615 497
rect 561 451 571 485
rect 605 451 615 485
rect 561 413 615 451
rect 645 413 711 497
rect 741 485 802 497
rect 741 451 760 485
rect 794 451 802 485
rect 741 413 802 451
rect 856 485 908 497
rect 856 451 864 485
rect 898 451 908 485
rect 465 369 515 413
rect 856 297 908 451
rect 938 471 992 497
rect 938 437 948 471
rect 982 437 992 471
rect 938 368 992 437
rect 938 334 948 368
rect 982 334 992 368
rect 938 297 992 334
rect 1022 489 1088 497
rect 1022 455 1038 489
rect 1072 455 1088 489
rect 1022 421 1088 455
rect 1022 387 1038 421
rect 1072 387 1088 421
rect 1022 297 1088 387
rect 1118 477 1179 497
rect 1118 443 1131 477
rect 1165 443 1179 477
rect 1118 297 1179 443
rect 1209 475 1261 497
rect 1209 441 1219 475
rect 1253 441 1261 475
rect 1209 384 1261 441
rect 1209 350 1219 384
rect 1253 350 1261 384
rect 1209 297 1261 350
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 85 341 119
rect 391 55 425 89
rect 867 131 901 165
rect 579 73 613 107
rect 763 72 797 106
rect 867 63 901 97
rect 1035 55 1069 89
rect 1135 55 1169 89
rect 1219 59 1253 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 449 341 483
rect 307 381 341 415
rect 391 451 425 485
rect 391 383 425 417
rect 571 451 605 485
rect 760 451 794 485
rect 864 451 898 485
rect 948 437 982 471
rect 948 334 982 368
rect 1038 455 1072 489
rect 1038 387 1072 421
rect 1131 443 1165 477
rect 1219 441 1253 475
rect 1219 350 1253 384
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 435 497 465 523
rect 531 497 561 523
rect 615 497 645 523
rect 711 497 741 523
rect 908 497 938 523
rect 992 497 1022 523
rect 1088 497 1118 523
rect 1179 497 1209 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 280 76 318
rect 21 264 76 280
rect 163 274 193 363
rect 21 230 32 264
rect 66 230 76 264
rect 21 214 76 230
rect 118 264 193 274
rect 118 230 134 264
rect 168 230 193 264
rect 351 241 381 369
rect 118 220 193 230
rect 46 176 76 214
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 298 225 381 241
rect 298 191 308 225
rect 342 191 381 225
rect 435 219 465 369
rect 531 337 561 413
rect 615 375 645 413
rect 507 321 561 337
rect 603 365 669 375
rect 603 331 619 365
rect 653 331 669 365
rect 603 321 669 331
rect 711 373 741 413
rect 711 357 812 373
rect 711 323 768 357
rect 802 323 812 357
rect 507 287 517 321
rect 551 287 561 321
rect 711 307 812 323
rect 507 279 561 287
rect 507 271 658 279
rect 531 249 658 271
rect 298 175 381 191
rect 351 131 381 175
rect 423 203 477 219
rect 423 169 433 203
rect 467 169 477 203
rect 423 153 477 169
rect 519 197 586 207
rect 519 163 536 197
rect 570 163 586 197
rect 519 153 586 163
rect 435 131 465 153
rect 530 119 560 153
rect 628 119 658 249
rect 723 131 753 307
rect 908 260 938 297
rect 992 265 1022 297
rect 1088 265 1118 297
rect 1179 265 1209 297
rect 908 259 941 260
rect 796 249 941 259
rect 796 215 812 249
rect 846 215 941 249
rect 796 205 941 215
rect 911 177 941 205
rect 983 249 1037 265
rect 983 215 993 249
rect 1027 215 1037 249
rect 983 199 1037 215
rect 1079 249 1209 265
rect 1079 215 1089 249
rect 1123 215 1209 249
rect 1079 199 1209 215
rect 995 177 1025 199
rect 1095 177 1125 199
rect 1179 177 1209 199
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 435 21 465 47
rect 530 21 560 47
rect 628 21 658 47
rect 723 21 753 47
rect 911 21 941 47
rect 995 21 1025 47
rect 1095 21 1125 47
rect 1179 21 1209 47
<< polycont >>
rect 32 230 66 264
rect 134 230 168 264
rect 308 191 342 225
rect 619 331 653 365
rect 768 323 802 357
rect 517 287 551 321
rect 433 169 467 203
rect 536 163 570 197
rect 812 215 846 249
rect 993 215 1027 249
rect 1089 215 1123 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 391 485 454 527
rect 760 485 822 527
rect 237 443 248 477
rect 203 409 248 443
rect 69 375 156 393
rect 35 359 156 375
rect 17 264 66 325
rect 17 230 32 264
rect 17 197 66 230
rect 122 323 156 359
rect 122 280 156 289
rect 237 391 248 409
rect 203 357 214 375
rect 203 337 248 357
rect 291 449 307 483
rect 341 449 357 483
rect 291 415 357 449
rect 291 381 307 415
rect 341 381 357 415
rect 122 264 168 280
rect 122 230 134 264
rect 122 214 168 230
rect 122 161 156 214
rect 35 127 156 161
rect 35 119 69 127
rect 203 119 237 337
rect 291 333 357 381
rect 425 451 454 485
rect 555 451 571 485
rect 605 451 721 485
rect 391 417 454 451
rect 425 383 454 417
rect 391 367 454 383
rect 494 391 551 401
rect 528 357 551 391
rect 291 299 428 333
rect 292 225 358 265
rect 292 191 308 225
rect 342 191 358 225
rect 392 219 428 299
rect 494 321 551 357
rect 494 287 517 321
rect 494 271 551 287
rect 585 365 653 399
rect 585 331 619 365
rect 585 323 653 331
rect 585 289 586 323
rect 620 289 653 323
rect 585 283 653 289
rect 585 229 619 283
rect 687 265 721 451
rect 794 451 822 485
rect 760 427 822 451
rect 856 485 912 527
rect 856 451 864 485
rect 898 451 912 485
rect 856 427 912 451
rect 946 471 984 493
rect 946 437 948 471
rect 982 437 984 471
rect 946 373 984 437
rect 1018 489 1092 527
rect 1018 455 1038 489
rect 1072 455 1092 489
rect 1018 421 1092 455
rect 1018 387 1038 421
rect 1072 387 1092 421
rect 1018 375 1092 387
rect 1131 477 1185 493
rect 1165 443 1185 477
rect 1131 375 1185 443
rect 764 368 984 373
rect 764 357 948 368
rect 764 323 768 357
rect 802 334 948 357
rect 982 341 984 368
rect 982 334 1117 341
rect 802 323 1117 334
rect 764 307 1117 323
rect 1083 265 1117 307
rect 1151 300 1185 375
rect 1219 475 1271 527
rect 1253 441 1271 475
rect 1219 384 1271 441
rect 1253 350 1271 384
rect 1219 334 1271 350
rect 1151 285 1271 300
rect 1152 283 1271 285
rect 1153 282 1271 283
rect 1155 277 1271 282
rect 687 249 862 265
rect 392 203 468 219
rect 392 169 433 203
rect 467 169 468 203
rect 392 157 468 169
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 203 69 237 85
rect 307 153 468 157
rect 535 197 619 229
rect 535 163 536 197
rect 570 163 619 197
rect 307 123 428 153
rect 535 141 619 163
rect 666 215 812 249
rect 846 215 862 249
rect 666 205 862 215
rect 896 249 1034 265
rect 896 215 993 249
rect 1027 215 1034 249
rect 307 119 341 123
rect 666 107 700 205
rect 896 199 1034 215
rect 1070 249 1123 265
rect 1070 215 1089 249
rect 1070 199 1123 215
rect 1083 165 1117 199
rect 1157 178 1271 277
rect 1154 173 1271 178
rect 307 69 341 85
rect 103 17 169 59
rect 375 55 391 89
rect 425 55 441 89
rect 562 73 579 107
rect 613 73 700 107
rect 848 131 867 165
rect 901 131 1117 165
rect 1151 153 1271 173
rect 375 17 441 55
rect 747 72 763 106
rect 797 72 814 106
rect 747 17 814 72
rect 848 97 918 131
rect 1151 97 1185 153
rect 848 63 867 97
rect 901 63 918 97
rect 848 51 918 63
rect 1019 89 1085 97
rect 1019 55 1035 89
rect 1069 55 1085 89
rect 1019 17 1085 55
rect 1119 89 1185 97
rect 1119 55 1135 89
rect 1169 55 1185 89
rect 1119 51 1185 55
rect 1219 93 1271 119
rect 1253 59 1271 93
rect 1219 17 1271 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 122 289 156 323
rect 214 375 237 391
rect 237 375 248 391
rect 214 357 248 375
rect 494 357 528 391
rect 586 289 620 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 482 391 540 397
rect 482 388 494 391
rect 248 360 494 388
rect 248 357 260 360
rect 202 351 260 357
rect 482 357 494 360
rect 528 357 540 391
rect 482 351 540 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 574 323 632 329
rect 574 320 586 323
rect 156 292 586 320
rect 156 289 168 292
rect 110 283 168 289
rect 574 289 586 292
rect 620 289 632 323
rect 574 283 632 289
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel locali s 954 221 988 255 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1138 425 1172 459 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1227 153 1261 187 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1227 221 1261 255 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 310 221 344 255 0 FreeSans 200 0 0 0 D
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew clock input
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
flabel metal1 s 46 544 46 544 0 FreeSans 200 0 0 0 VPWR
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel nwell s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
flabel nwell s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel pwell s 47 0 47 0 0 FreeSans 200 0 0 0 VNB
flabel pwell s 47 0 47 0 0 FreeSans 200 0 0 0 VNB
rlabel comment s 0 0 0 0 4 dlrtn_2
rlabel metal1 s 0 -48 1288 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1288 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_END 2763190
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2751784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
