magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< mvpmos >>
tri 3574 3903 3594 3923 sw
tri 6654 3903 6674 3923 se
rect 3574 3793 6674 3903
tri 3574 3773 3594 3793 nw
tri 6654 3773 6674 3793 ne
tri 6816 3903 6836 3923 sw
tri 9896 3903 9916 3923 se
rect 6816 3793 9916 3903
tri 6816 3773 6836 3793 nw
tri 9896 3773 9916 3793 ne
tri 10058 3903 10078 3923 sw
tri 13138 3903 13158 3923 se
rect 10058 3793 13158 3903
tri 10058 3773 10078 3793 nw
tri 13138 3773 13158 3793 ne
tri 13300 3903 13320 3923 sw
tri 16380 3903 16400 3923 se
rect 13300 3793 16400 3903
tri 13300 3773 13320 3793 nw
tri 16380 3773 16400 3793 ne
tri 16542 3903 16562 3923 sw
tri 19622 3903 19642 3923 se
rect 16542 3793 19642 3903
tri 16542 3773 16562 3793 nw
tri 19622 3773 19642 3793 ne
tri 19784 3903 19804 3923 sw
tri 22864 3903 22884 3923 se
rect 19784 3793 22884 3903
tri 19784 3773 19804 3793 nw
tri 22864 3773 22884 3793 ne
tri 3574 3491 3594 3511 sw
tri 6654 3491 6674 3511 se
rect 3574 3381 6674 3491
tri 3574 3361 3594 3381 nw
tri 6654 3361 6674 3381 ne
tri 6816 3491 6836 3511 sw
tri 9896 3491 9916 3511 se
rect 6816 3381 9916 3491
tri 6816 3361 6836 3381 nw
tri 9896 3361 9916 3381 ne
tri 10058 3491 10078 3511 sw
tri 13138 3491 13158 3511 se
rect 10058 3381 13158 3491
tri 10058 3361 10078 3381 nw
tri 13138 3361 13158 3381 ne
tri 13300 3491 13320 3511 sw
tri 16380 3491 16400 3511 se
rect 13300 3381 16400 3491
tri 13300 3361 13320 3381 nw
tri 16380 3361 16400 3381 ne
tri 16542 3491 16562 3511 sw
tri 19622 3491 19642 3511 se
rect 16542 3381 19642 3491
tri 16542 3361 16562 3381 nw
tri 19622 3361 19642 3381 ne
tri 19784 3491 19804 3511 sw
tri 22864 3491 22884 3511 se
rect 19784 3381 22884 3491
tri 19784 3361 19804 3381 nw
tri 22864 3361 22884 3381 ne
<< poly >>
rect 23025 7319 23075 7352
rect 23025 7285 23041 7319
rect 23025 7252 23075 7285
rect 25115 7319 25165 7352
rect 25149 7285 25165 7319
rect 25115 7252 25165 7285
rect 23016 7093 23066 7126
rect 23016 7059 23032 7093
rect 23016 7026 23066 7059
rect 25106 7093 25156 7126
rect 25140 7059 25156 7093
rect 25106 7026 25156 7059
<< polycont >>
rect 23041 7285 23075 7319
rect 25115 7285 25149 7319
rect 23032 7059 23066 7093
rect 25106 7059 25140 7093
<< npolyres >>
rect 23075 7252 25115 7352
rect 23066 7026 25106 7126
<< locali >>
rect 23041 7320 23075 7335
rect 23071 7319 23109 7320
rect 23075 7286 23109 7319
rect 23041 7269 23075 7285
rect 23053 7093 23066 7109
rect 23019 7059 23032 7083
rect 23019 7045 23066 7059
rect 23053 7043 23066 7045
<< viali >>
rect 23037 7319 23071 7320
rect 23037 7286 23041 7319
rect 23041 7286 23071 7319
rect 23109 7286 23143 7320
rect 25115 7319 25221 7348
rect 25115 7285 25149 7319
rect 25149 7285 25221 7319
rect 25115 7242 25221 7285
rect 23019 7093 23053 7117
rect 23019 7083 23032 7093
rect 23032 7083 23053 7093
rect 23019 7011 23053 7045
rect 25106 7093 25212 7116
rect 25106 7059 25140 7093
rect 25140 7059 25212 7093
rect 25106 7010 25212 7059
<< metal1 >>
rect 777 16922 823 16974
tri 777 16920 779 16922 ne
rect 779 16920 823 16922
tri 1931 16708 1960 16737 ne
tri 199 16610 227 16638 ne
rect 227 16610 233 16638
tri 227 16604 233 16610 ne
rect 285 16610 291 16638
tri 291 16610 319 16638 nw
tri 285 16604 291 16610 nw
rect 1644 16561 1734 16610
tri 1644 16558 1647 16561 ne
rect 1647 16558 1734 16561
rect 1862 16558 1907 16610
tri 285 16492 319 16526 sw
tri 601 16492 607 16498 sw
rect 285 16434 313 16440
tri 313 16434 319 16440 nw
tri 285 16406 313 16434 nw
rect 601 16355 607 16492
tri 1835 16430 1839 16434 se
rect 1839 16430 1841 16434
rect 1964 16430 1969 16434
tri 1969 16430 1973 16434 sw
rect 1835 16391 1973 16430
tri 1830 16382 1839 16391 ne
rect 1839 16386 1973 16391
rect 1839 16382 1969 16386
tri 1969 16382 1973 16386 nw
tri 601 16349 607 16355 nw
tri 549 16185 555 16191 se
rect 549 16048 555 16185
tri 549 16042 555 16048 ne
tri 1009 15889 1025 15905 sw
rect 803 15883 1025 15889
rect 803 15831 804 15883
rect 856 15831 888 15883
rect 940 15831 972 15883
rect 1024 15831 1025 15883
rect 803 15804 1025 15831
rect 803 15752 804 15804
rect 856 15752 888 15804
rect 940 15752 972 15804
rect 1024 15752 1025 15804
rect 803 15725 1025 15752
rect 803 15673 804 15725
rect 856 15673 888 15725
rect 940 15673 972 15725
rect 1024 15673 1025 15725
rect 803 15646 1025 15673
rect 803 15594 804 15646
rect 856 15594 888 15646
rect 940 15594 972 15646
rect 1024 15594 1025 15646
rect 803 15588 1025 15594
tri 1009 15572 1025 15588 nw
tri 744 14613 778 14647 se
tri 744 14562 749 14567 ne
rect 749 14562 778 14567
rect 549 14425 555 14562
tri 749 14533 778 14562 ne
tri 549 14419 555 14425 ne
rect 932 12912 1002 13195
tri 549 12707 555 12713 se
rect 549 12568 555 12707
tri 549 12562 555 12568 ne
tri 876 8376 901 8401 ne
rect 901 8376 910 8401
rect 25109 7353 25227 7360
rect 23025 7277 23031 7329
rect 23083 7277 23097 7329
rect 23149 7277 23155 7329
rect 2671 7186 2692 7238
rect 25225 7237 25227 7353
rect 25109 7230 25227 7237
rect 23013 7122 23065 7129
rect 23013 7058 23065 7070
rect 23013 6999 23065 7006
rect 25100 7122 25221 7128
rect 25100 7006 25105 7122
rect 25100 6998 25221 7006
rect 6333 6480 6339 6532
rect 6391 6480 6405 6532
rect 6457 6480 6471 6532
rect 6523 6480 6537 6532
rect 6589 6480 6603 6532
rect 6655 6480 6668 6532
rect 6720 6480 6733 6532
rect 6785 6480 6798 6532
rect 6850 6480 6863 6532
rect 6915 6480 6928 6532
rect 6980 6480 6993 6532
rect 7045 6480 7058 6532
rect 7110 6480 7123 6532
rect 7175 6480 7188 6532
rect 7240 6480 7253 6532
rect 7305 6480 7318 6532
rect 7370 6480 7383 6532
rect 7435 6480 7448 6532
rect 7500 6480 7513 6532
rect 7565 6480 7578 6532
rect 7630 6480 7636 6532
rect 6333 6416 7636 6480
rect 6333 6364 6339 6416
rect 6391 6364 6405 6416
rect 6457 6364 6471 6416
rect 6523 6364 6537 6416
rect 6589 6364 6603 6416
rect 6655 6364 6668 6416
rect 6720 6364 6733 6416
rect 6785 6364 6798 6416
rect 6850 6364 6863 6416
rect 6915 6364 6928 6416
rect 6980 6364 6993 6416
rect 7045 6364 7058 6416
rect 7110 6364 7123 6416
rect 7175 6364 7188 6416
rect 7240 6364 7253 6416
rect 7305 6364 7318 6416
rect 7370 6364 7383 6416
rect 7435 6364 7448 6416
rect 7500 6364 7513 6416
rect 7565 6364 7578 6416
rect 7630 6364 7636 6416
rect 18353 6480 18359 6532
rect 18411 6480 18428 6532
rect 18480 6480 18497 6532
rect 18549 6480 18565 6532
rect 18617 6480 18633 6532
rect 18685 6480 18701 6532
rect 18753 6480 18769 6532
rect 18821 6480 18837 6532
rect 18889 6480 18905 6532
rect 18957 6480 18973 6532
rect 19025 6480 19041 6532
rect 19093 6480 19109 6532
rect 19161 6480 19177 6532
rect 19229 6480 19235 6532
rect 18353 6416 19235 6480
rect 18353 6364 18359 6416
rect 18411 6364 18428 6416
rect 18480 6364 18497 6416
rect 18549 6364 18565 6416
rect 18617 6364 18633 6416
rect 18685 6364 18701 6416
rect 18753 6364 18769 6416
rect 18821 6364 18837 6416
rect 18889 6364 18905 6416
rect 18957 6364 18973 6416
rect 19025 6364 19041 6416
rect 19093 6364 19109 6416
rect 19161 6364 19177 6416
rect 19229 6364 19235 6416
rect 20192 6480 20198 6532
rect 20250 6480 20267 6532
rect 20319 6480 20336 6532
rect 20388 6480 20404 6532
rect 20456 6480 20472 6532
rect 20524 6480 20540 6532
rect 20592 6480 20608 6532
rect 20660 6480 20676 6532
rect 20728 6480 20744 6532
rect 20796 6480 20812 6532
rect 20864 6480 20880 6532
rect 20932 6480 20948 6532
rect 21000 6480 21016 6532
rect 21068 6480 21074 6532
rect 20192 6416 21074 6480
rect 20192 6364 20198 6416
rect 20250 6364 20267 6416
rect 20319 6364 20336 6416
rect 20388 6364 20404 6416
rect 20456 6364 20472 6416
rect 20524 6364 20540 6416
rect 20592 6364 20608 6416
rect 20660 6364 20676 6416
rect 20728 6364 20744 6416
rect 20796 6364 20812 6416
rect 20864 6364 20880 6416
rect 20932 6364 20948 6416
rect 21000 6364 21016 6416
rect 21068 6364 21074 6416
rect 22975 6480 22981 6532
rect 23033 6480 23072 6532
rect 23124 6480 23130 6532
rect 22975 6416 23130 6480
rect 22975 6364 22981 6416
rect 23033 6364 23072 6416
rect 23124 6364 23130 6416
tri 23152 5777 23154 5779 se
rect 23154 5773 23270 5779
tri 23270 5777 23272 5779 sw
rect 23154 5587 23270 5593
rect 1753 5468 1936 5552
rect 8088 5498 8094 5550
rect 8146 5498 8158 5550
rect 8210 5498 8216 5550
rect 11308 5498 11314 5550
rect 11366 5498 11378 5550
rect 11430 5498 11436 5550
rect 14528 5498 14534 5550
rect 14586 5498 14598 5550
rect 14650 5498 14656 5550
rect 17748 5498 17754 5550
rect 17806 5498 17818 5550
rect 17870 5498 17876 5550
rect 20968 5498 20974 5550
rect 21026 5498 21038 5550
rect 21090 5498 21096 5550
rect 24188 5498 24194 5550
rect 24246 5498 24258 5550
rect 24310 5498 24316 5550
tri 26003 5439 26032 5468 ne
rect 26032 5439 26051 5468
tri 6114 5387 6121 5394 ne
rect 6121 5387 6127 5439
rect 6179 5387 6191 5439
rect 6243 5387 6249 5439
tri 6249 5387 6256 5394 nw
rect 25548 5393 25583 5439
tri 25548 5387 25554 5393 ne
rect 25554 5387 25583 5393
tri 25554 5364 25577 5387 ne
tri 3029 5358 3035 5364 se
rect 3035 5312 3041 5364
rect 3093 5312 3105 5364
rect 3157 5312 3163 5364
tri 3163 5358 3169 5364 sw
tri 3561 5358 3567 5364 se
rect 3567 5358 3695 5364
tri 3695 5358 3701 5364 sw
rect 25577 5323 25583 5387
rect 25699 5323 25705 5439
tri 26032 5420 26051 5439 ne
tri 25838 5284 25842 5288 se
rect 25842 5284 25958 5288
tri 2880 5280 2884 5284 sw
tri 25836 5282 25838 5284 se
rect 25838 5282 25958 5284
rect 2880 5248 2896 5280
rect 2880 5242 2890 5248
tri 2890 5242 2896 5248 nw
rect 2435 5190 2441 5242
rect 2493 5190 2505 5242
rect 2557 5232 2563 5242
rect 2880 5237 2885 5242
tri 2885 5237 2890 5242 nw
tri 2563 5232 2568 5237 sw
tri 2880 5232 2885 5237 nw
rect 2557 5217 2568 5232
tri 2568 5217 2583 5232 sw
rect 2557 5201 2699 5217
tri 2699 5201 2715 5217 sw
tri 2896 5201 2912 5217 se
rect 2912 5201 16270 5217
rect 2557 5190 16270 5201
rect 2435 5185 16270 5190
tri 2659 5169 2675 5185 ne
rect 2675 5169 2934 5185
tri 2934 5169 2950 5185 nw
tri 16244 5169 16260 5185 ne
rect 16260 5169 16270 5185
tri 16260 5166 16263 5169 ne
rect 16263 5166 16270 5169
tri 16263 5165 16264 5166 ne
rect 16264 5165 16270 5166
rect 16322 5165 16337 5217
rect 16389 5165 16404 5217
rect 16456 5165 16470 5217
rect 16522 5165 16528 5217
rect 23347 5166 23353 5282
rect 23469 5266 25842 5282
rect 23469 5214 24798 5266
rect 24850 5214 24862 5266
rect 24914 5214 25842 5266
rect 23469 5197 25842 5214
rect 23469 5166 23475 5197
tri 23475 5166 23506 5197 nw
tri 25805 5166 25836 5197 ne
rect 25836 5166 25842 5197
tri 25836 5165 25837 5166 ne
rect 25837 5165 25958 5166
tri 25837 5160 25842 5165 ne
rect 25842 5160 25958 5165
rect 2508 5103 2514 5155
rect 2566 5103 2578 5155
rect 2630 5131 2636 5155
tri 2636 5131 2660 5155 sw
tri 2948 5131 2972 5155 se
rect 2972 5131 9390 5155
rect 2630 5124 9390 5131
tri 9390 5124 9421 5155 sw
rect 2630 5123 9421 5124
rect 2630 5103 2975 5123
tri 2975 5103 2995 5123 nw
tri 9337 5103 9357 5123 ne
rect 9357 5103 9421 5123
tri 9357 5093 9367 5103 ne
rect 9367 5093 9421 5103
tri 8390 5087 8396 5093 se
rect 8396 5087 8524 5093
tri 8524 5087 8530 5093 sw
tri 9367 5089 9371 5093 ne
rect 8390 5085 8530 5087
tri 8530 5085 8532 5087 sw
rect 8390 5049 8532 5085
rect 8390 5047 8530 5049
tri 8530 5047 8532 5049 nw
tri 8390 5041 8396 5047 ne
rect 8396 5041 8524 5047
tri 8524 5041 8530 5047 nw
rect 6274 4966 6280 5018
rect 6332 4966 6344 5018
rect 6396 4966 7638 5018
rect 7690 4966 7702 5018
rect 7754 4966 7760 5018
rect 9371 4966 9421 5093
tri 11610 5087 11616 5093 se
rect 11616 5087 11745 5093
tri 11745 5087 11751 5093 sw
rect 11610 5086 11751 5087
tri 11751 5086 11752 5087 sw
rect 11610 5048 11752 5086
rect 11610 5047 11751 5048
tri 11751 5047 11752 5048 nw
rect 18050 5047 18190 5093
tri 11610 5041 11616 5047 ne
rect 11616 5041 11745 5047
tri 11745 5041 11751 5047 nw
tri 14830 5041 14836 5047 ne
rect 14836 5041 14964 5047
tri 14964 5041 14970 5047 nw
tri 18050 5041 18056 5047 ne
rect 18056 5041 18184 5047
tri 18184 5041 18190 5047 nw
rect 21270 5047 21410 5093
tri 21270 5041 21276 5047 ne
rect 21276 5041 21404 5047
tri 21404 5041 21410 5047 nw
rect 24490 5047 24630 5093
tri 24490 5041 24496 5047 ne
rect 24496 5041 24624 5047
tri 24624 5041 24630 5047 nw
tri 9421 4966 9431 4976 sw
rect 9371 4940 9431 4966
tri 9431 4940 9457 4966 sw
rect 5423 4888 5429 4940
rect 5481 4888 5507 4940
rect 5559 4888 5585 4940
rect 5637 4888 5643 4940
tri 7830 4937 7833 4940 se
rect 7833 4937 7839 4940
rect 7830 4891 7839 4937
tri 7830 4888 7833 4891 ne
rect 7833 4888 7839 4891
rect 7891 4888 7908 4940
rect 7960 4888 7976 4940
rect 8028 4937 8034 4940
tri 8034 4937 8037 4940 sw
rect 8028 4891 8037 4937
rect 9371 4937 9457 4940
tri 9457 4937 9460 4940 sw
tri 13441 4937 13444 4940 se
rect 13444 4937 13450 4940
rect 9371 4923 9470 4937
tri 9371 4891 9403 4923 ne
rect 9403 4891 9470 4923
rect 9489 4897 9521 4929
rect 13441 4891 13450 4937
rect 8028 4888 8034 4891
tri 8034 4888 8037 4891 nw
tri 13441 4888 13444 4891 ne
rect 13444 4888 13450 4891
rect 13502 4888 13519 4940
rect 13571 4888 13587 4940
rect 13639 4937 13645 4940
tri 13645 4937 13648 4940 sw
rect 13639 4891 13648 4937
rect 13639 4888 13645 4891
tri 13645 4888 13648 4891 nw
tri 16261 4937 16264 4940 se
rect 16264 4937 16270 4940
rect 16261 4891 16270 4937
tri 16261 4888 16264 4891 ne
rect 16264 4888 16270 4891
rect 16322 4888 16337 4940
rect 16389 4888 16404 4940
rect 16456 4888 16470 4940
rect 16522 4937 16528 4940
tri 16528 4937 16531 4940 sw
rect 16522 4891 16531 4937
rect 16522 4888 16528 4891
tri 16528 4888 16531 4891 nw
tri 19510 4937 19513 4940 se
rect 19513 4937 19519 4940
rect 19510 4891 19519 4937
tri 19510 4888 19513 4891 ne
rect 19513 4888 19519 4891
rect 19571 4888 19588 4940
rect 19640 4888 19656 4940
rect 19708 4937 19714 4940
tri 19714 4937 19717 4940 sw
rect 19708 4891 19717 4937
rect 19708 4888 19714 4891
tri 19714 4888 19717 4891 nw
tri 22904 4937 22907 4940 se
rect 22907 4937 22913 4940
rect 22904 4891 22913 4937
tri 22904 4888 22907 4891 ne
rect 22907 4888 22913 4891
rect 22965 4888 22982 4940
rect 23034 4888 23050 4940
rect 23102 4937 23108 4940
tri 23108 4937 23111 4940 sw
rect 23102 4891 23111 4937
rect 23102 4888 23108 4891
tri 23108 4888 23111 4891 nw
rect 2680 4734 2686 4786
rect 2738 4734 2750 4786
rect 2802 4784 2808 4786
tri 2808 4784 2810 4786 sw
rect 2802 4781 2810 4784
tri 2810 4781 2813 4784 sw
tri 8393 4781 8396 4784 se
rect 8396 4781 8524 4784
tri 8524 4781 8527 4784 sw
rect 2802 4735 3298 4781
rect 8393 4735 8527 4781
rect 2802 4734 2808 4735
tri 2808 4734 2809 4735 nw
tri 8393 4734 8394 4735 ne
rect 8394 4734 8524 4735
tri 8394 4732 8396 4734 ne
rect 8396 4732 8524 4734
tri 8524 4732 8527 4735 nw
tri 11610 4778 11616 4784 se
rect 11616 4778 11745 4784
tri 11745 4778 11751 4784 sw
tri 14833 4781 14836 4784 se
rect 14836 4781 14964 4784
tri 14964 4781 14967 4784 sw
rect 11610 4777 11751 4778
tri 11751 4777 11752 4778 sw
rect 11610 4739 11752 4777
rect 11610 4738 11751 4739
tri 11751 4738 11752 4739 nw
tri 11610 4732 11616 4738 ne
rect 11616 4732 11745 4738
tri 11745 4732 11751 4738 nw
rect 14833 4735 14967 4781
tri 14833 4732 14836 4735 ne
rect 14836 4732 14964 4735
tri 14964 4732 14967 4735 nw
tri 18053 4781 18056 4784 se
rect 18056 4781 18184 4784
tri 18184 4781 18187 4784 sw
rect 18053 4735 18187 4781
tri 18053 4732 18056 4735 ne
rect 18056 4732 18184 4735
tri 18184 4732 18187 4735 nw
tri 21273 4781 21276 4784 se
rect 21276 4781 21404 4784
tri 21404 4781 21407 4784 sw
rect 21273 4735 21407 4781
tri 21273 4732 21276 4735 ne
rect 21276 4732 21404 4735
tri 21404 4732 21407 4735 nw
tri 24493 4781 24496 4784 se
rect 24496 4781 24624 4784
tri 24624 4781 24627 4784 sw
rect 24493 4735 24627 4781
tri 24493 4732 24496 4735 ne
rect 24496 4732 24624 4735
tri 24624 4732 24627 4735 nw
tri 3058 4700 3064 4706 se
rect 3064 4700 3192 4706
tri 3192 4700 3198 4706 sw
rect 1625 4681 2775 4686
tri 2775 4681 2780 4686 sw
rect 1625 4660 2780 4681
tri 2780 4660 2801 4681 sw
rect 1625 4654 2801 4660
tri 2752 4626 2780 4654 ne
rect 2780 4626 2801 4654
tri 2801 4626 2835 4660 sw
tri 25702 4626 25736 4660 se
rect 25736 4626 25742 4660
tri 2780 4595 2811 4626 ne
rect 2811 4595 22913 4626
rect 1625 4594 2767 4595
tri 2767 4594 2768 4595 sw
tri 2811 4594 2812 4595 ne
rect 2812 4594 22913 4595
rect 1625 4574 2768 4594
tri 2768 4574 2788 4594 sw
tri 22887 4574 22907 4594 ne
rect 22907 4574 22913 4594
rect 22965 4574 22982 4626
rect 23034 4574 23050 4626
rect 23102 4594 23560 4626
tri 25692 4616 25702 4626 se
rect 25702 4616 25742 4626
rect 23102 4574 23108 4594
tri 23108 4574 23128 4594 nw
rect 1625 4566 2788 4574
tri 2788 4566 2796 4574 sw
rect 1625 4563 19519 4566
tri 2744 4534 2773 4563 ne
rect 2773 4534 19519 4563
tri 19493 4514 19513 4534 ne
rect 19513 4514 19519 4534
rect 19571 4514 19588 4566
rect 19640 4514 19656 4566
rect 19708 4541 22869 4566
tri 22869 4541 22894 4566 sw
rect 19708 4534 23464 4541
rect 19708 4514 19714 4534
tri 19714 4514 19734 4534 nw
tri 22827 4514 22847 4534 ne
rect 22847 4514 23464 4534
tri 22847 4509 22852 4514 ne
rect 22852 4509 23464 4514
tri 23377 4506 23380 4509 ne
rect 23380 4506 23464 4509
rect 2762 4474 7839 4506
tri 7813 4454 7833 4474 ne
rect 7833 4454 7839 4474
rect 7891 4454 7908 4506
rect 7960 4454 7976 4506
rect 8028 4454 8034 4506
rect 8086 4454 8092 4506
rect 8144 4454 8156 4506
rect 8208 4454 8698 4506
rect 8750 4454 8762 4506
rect 8814 4454 11918 4506
rect 11970 4454 11982 4506
rect 12034 4454 13219 4506
rect 13271 4454 13283 4506
rect 13335 4473 13787 4506
rect 13335 4454 13395 4473
tri 13395 4454 13414 4473 nw
tri 13660 4454 13679 4473 ne
rect 13679 4454 13787 4473
rect 13839 4454 13851 4506
rect 13903 4454 15138 4506
rect 15190 4454 15202 4506
rect 15254 4454 18358 4506
rect 18410 4454 18422 4506
rect 18474 4454 19299 4506
rect 19351 4454 19363 4506
rect 19415 4500 19457 4506
tri 19457 4500 19463 4506 sw
tri 19752 4500 19758 4506 se
rect 19758 4500 19867 4506
rect 19415 4485 19463 4500
tri 19463 4485 19478 4500 sw
tri 19737 4485 19752 4500 se
rect 19752 4485 19867 4500
rect 19415 4454 19867 4485
rect 19919 4454 19931 4506
rect 19983 4454 21578 4506
rect 21630 4454 21642 4506
rect 21694 4454 22636 4506
rect 22688 4454 22700 4506
rect 22752 4454 22758 4506
tri 23380 4500 23386 4506 ne
rect 23386 4500 23464 4506
rect 23657 4500 23663 4616
rect 23779 4544 25742 4616
rect 25858 4544 25864 4660
rect 23779 4500 23785 4544
tri 23785 4500 23829 4544 nw
tri 23386 4474 23412 4500 ne
tri 13424 4424 13444 4444 se
rect 13444 4424 13450 4444
rect 3044 4392 13450 4424
rect 13502 4392 13519 4444
rect 13571 4392 13587 4444
rect 13639 4424 13645 4444
tri 13645 4424 13665 4444 sw
rect 13639 4392 23368 4424
rect 22920 3831 22972 3914
tri 3454 3493 3466 3505 se
rect 2844 2470 3047 2476
rect 2896 2418 2995 2470
rect 2844 2406 3047 2418
rect 2896 2354 2995 2406
rect 2844 2348 3047 2354
rect 2326 1758 2896 1764
rect 2378 1706 2844 1758
rect 2326 1694 2896 1706
rect 2378 1642 2844 1694
rect 2326 1636 2896 1642
tri 2996 1344 2997 1345 ne
rect 2997 1344 2999 1345
rect 23412 1135 23464 4500
rect 23654 2860 23734 2907
tri 23624 2811 23654 2841 se
rect 23654 2811 23734 2858
tri 23734 2811 23765 2842 sw
rect 23602 2731 23811 2811
rect 23813 2731 23860 2811
rect 23602 1306 23687 2731
tri 23687 2675 23743 2731 nw
tri 23602 1292 23616 1306 ne
rect 23616 1292 23687 1306
tri 23687 1292 23744 1349 sw
tri 23616 1221 23687 1292 ne
rect 23687 1280 23789 1292
rect 23687 1228 23720 1280
rect 23772 1228 23789 1280
rect 23687 1221 23789 1228
tri 23687 1204 23704 1221 ne
rect 23704 1216 23789 1221
rect 23704 1164 23720 1216
rect 23772 1164 23789 1216
rect 23704 1152 23789 1164
rect 23704 1100 23720 1152
rect 23772 1100 23789 1152
rect 23704 1094 23789 1100
tri 2378 993 2408 1023 sw
rect 2451 947 2491 993
tri 2294 915 2322 943 sw
tri 6615 861 6617 863 ne
rect 6617 861 6650 863
tri 2210 831 2240 861 sw
tri 6617 831 6647 861 ne
rect 6647 831 6650 861
tri 6647 828 6650 831 ne
tri 4719 821 4725 827 se
rect 4725 821 4728 827
tri 2126 775 2131 780 sw
rect 4719 775 4728 821
tri 4937 821 4943 827 se
rect 4943 821 4946 827
rect 4937 775 4946 821
rect 5068 823 5071 827
tri 5071 823 5075 827 sw
rect 5068 821 5075 823
tri 5075 821 5077 823 sw
rect 5068 775 5077 821
tri 6412 821 6414 823 sw
rect 6412 775 6414 821
rect 2126 773 2131 775
tri 2131 773 2133 775 sw
tri 6412 773 6414 775 nw
rect 2126 749 2133 773
tri 2133 749 2157 773 sw
rect 2126 748 2157 749
tri 2157 748 2158 749 sw
tri 3837 748 3838 749 sw
rect 2844 696 2850 748
rect 2902 696 2914 748
rect 2966 696 2972 748
rect 3837 742 3838 748
tri 3838 742 3844 748 sw
rect 3837 728 3844 742
rect 6837 699 6889 704
tri 2042 667 2069 694 sw
tri 1958 584 1987 613 sw
tri 1874 517 1879 522 sw
rect 1874 501 1879 517
tri 1879 501 1895 517 sw
tri 3349 501 3365 517 se
rect 3365 501 3370 517
rect 1874 500 1895 501
tri 1895 500 1896 501 sw
tri 3348 500 3349 501 se
rect 3349 500 3370 501
tri 14206 500 14207 501 se
rect 14207 500 23551 501
rect 1874 490 1896 500
tri 1896 490 1906 500 sw
tri 3338 490 3348 500 se
rect 3348 490 3370 500
tri 3337 489 3338 490 se
rect 3338 489 3370 490
tri 9211 497 9214 500 se
rect 9214 497 13486 500
tri 13486 497 13489 500 sw
rect 9211 451 13489 497
tri 9211 449 9213 451 ne
rect 9213 449 13486 451
tri 3528 446 3531 449 se
tri 3351 426 3363 438 ne
tri 1790 397 1806 413 sw
rect 3659 397 3660 449
tri 9213 448 9214 449 ne
rect 9214 448 13486 449
tri 13486 448 13489 451 nw
tri 14204 498 14206 500 se
rect 14206 498 23551 500
tri 23551 498 23554 501 sw
rect 14204 497 23554 498
tri 23554 497 23555 498 sw
rect 14204 452 23555 497
tri 14204 449 14207 452 ne
rect 14207 449 23552 452
tri 23552 449 23555 452 nw
tri 23832 449 23840 457 se
tri 23831 448 23832 449 se
rect 23832 448 23840 449
tri 23829 446 23831 448 se
rect 23831 446 23840 448
tri 3846 443 3849 446 sw
tri 4940 443 4943 446 se
rect 3846 397 3852 443
rect 4937 397 4943 443
rect 1790 394 1806 397
tri 1806 394 1809 397 sw
tri 3846 394 3849 397 nw
tri 4940 394 4943 397 ne
tri 5071 443 5074 446 sw
tri 23826 443 23829 446 se
rect 23829 443 23840 446
rect 5071 397 5077 443
tri 23803 420 23826 443 se
rect 23826 420 23840 443
tri 5071 394 5074 397 nw
rect 1790 379 1809 394
tri 1809 379 1824 394 sw
tri 23812 361 23825 374 ne
rect 23825 361 23840 374
tri 4722 358 4725 361 se
rect 3670 312 3676 358
rect 4719 312 4725 358
rect 3670 309 3673 312
tri 3673 309 3676 312 nw
tri 4722 309 4725 312 ne
tri 4853 358 4856 361 sw
tri 6820 358 6823 361 se
rect 4853 312 4859 358
rect 6820 312 6823 358
tri 23825 346 23840 361 ne
tri 4853 309 4856 312 nw
tri 6820 309 6823 312 ne
tri 9211 341 9214 344 se
rect 9214 341 13486 344
tri 13486 341 13489 344 sw
tri 3670 306 3673 309 nw
rect 9211 295 13489 341
tri 9211 292 9214 295 ne
rect 9214 292 13486 295
tri 13486 292 13489 295 nw
tri 13617 341 13620 344 se
rect 13620 341 22965 344
tri 22965 341 22968 344 sw
rect 13617 295 22968 341
tri 13617 292 13620 295 ne
rect 13620 292 22965 295
tri 22965 292 22968 295 nw
tri 23821 273 23840 292 se
tri 6011 271 6013 273 se
rect 6013 271 6143 273
tri 6143 271 6145 273 sw
tri 23819 271 23821 273 se
rect 23821 271 23840 273
tri 23812 264 23819 271 se
rect 23819 264 23840 271
tri 6638 218 6654 234 se
tri 6609 189 6638 218 se
rect 6638 189 6654 218
tri 23811 189 23840 218 ne
tri 6608 188 6609 189 se
rect 6609 188 6654 189
tri 9211 185 9214 188 se
rect 9214 185 13486 188
tri 13486 185 13489 188 sw
rect 9211 139 13489 185
tri 9211 136 9214 139 ne
rect 9214 136 13486 139
tri 13486 136 13489 139 nw
tri 13617 185 13620 188 se
rect 13620 185 22965 188
tri 22965 185 22968 188 sw
rect 13617 139 22968 185
tri 13617 136 13620 139 ne
rect 13620 136 22965 139
tri 22965 136 22968 139 nw
tri 23813 108 23840 135 se
tri 24034 95 24037 98 se
rect 24037 95 24912 98
tri 24912 95 24915 98 sw
tri 23811 58 23815 62 ne
rect 23815 58 23840 62
tri 3140 55 3143 58 se
rect 3143 55 3145 58
rect 3140 9 3145 55
tri 3140 6 3143 9 ne
rect 3143 6 3145 9
rect 7724 55 7726 58
tri 7726 55 7729 58 sw
rect 7724 9 7729 55
tri 23815 46 23827 58 ne
rect 23827 46 23840 58
rect 24034 49 24915 95
tri 24034 46 24037 49 ne
rect 24037 46 24912 49
tri 24912 46 24915 49 nw
tri 23827 33 23840 46 ne
rect 7724 6 7726 9
tri 7726 6 7729 9 nw
tri 9211 29 9214 32 se
rect 9214 29 23571 32
tri 23571 29 23574 32 sw
rect 9211 -17 23574 29
tri 9211 -20 9214 -17 ne
rect 9214 -20 23571 -17
tri 23571 -20 23574 -17 nw
tri 23839 -20 23840 -19 se
tri 2840 -24 2844 -20 se
rect 2844 -24 2850 -20
rect 2840 -68 2850 -24
tri 2840 -72 2844 -68 ne
rect 2844 -72 2850 -68
rect 2902 -72 2914 -20
rect 2966 -22 2974 -20
tri 2974 -22 2976 -20 sw
rect 2966 -68 2976 -22
tri 23811 -48 23839 -20 se
rect 23839 -48 23840 -20
rect 2966 -72 2972 -68
tri 2972 -72 2976 -68 nw
tri 3140 -101 3143 -98 se
rect 3143 -101 3145 -98
rect 3140 -147 3145 -101
tri 3140 -150 3143 -147 ne
rect 3143 -150 3145 -147
rect 7724 -101 7726 -98
tri 7726 -101 7729 -98 sw
rect 7724 -147 7729 -101
rect 7724 -150 7726 -147
tri 7726 -150 7729 -147 nw
tri 9211 -127 9214 -124 se
rect 9214 -127 13486 -124
tri 13486 -127 13489 -124 sw
rect 9211 -173 13489 -127
tri 9211 -176 9214 -173 ne
rect 9214 -176 13486 -173
tri 13486 -176 13489 -173 nw
tri 13617 -127 13620 -124 se
rect 13620 -127 22965 -124
tri 22965 -127 22968 -124 sw
rect 13617 -173 22968 -127
tri 13617 -176 13620 -173 ne
rect 13620 -176 22965 -173
tri 22965 -176 22968 -173 nw
rect 1599 -420 1830 -249
rect 2157 -481 23860 -472
rect 2157 -533 2163 -481
rect 2215 -533 2227 -481
rect 2279 -533 23674 -481
rect 23726 -533 23738 -481
rect 23790 -533 23802 -481
rect 23854 -533 23860 -481
rect 2157 -542 23860 -533
rect 13714 -1522 13720 -1470
rect 13772 -1522 13788 -1470
rect 13840 -1522 13856 -1470
rect 13908 -1522 13924 -1470
rect 13976 -1522 13992 -1470
rect 14044 -1522 14060 -1470
rect 14112 -1522 14128 -1470
rect 14180 -1522 14196 -1470
rect 14248 -1522 14264 -1470
rect 14316 -1522 14332 -1470
rect 14384 -1522 14400 -1470
rect 14452 -1522 14468 -1470
rect 14520 -1522 14536 -1470
rect 14588 -1522 14594 -1470
rect 18349 -1522 18355 -1470
rect 18407 -1522 18423 -1470
rect 18475 -1522 18491 -1470
rect 18543 -1522 18559 -1470
rect 18611 -1522 18627 -1470
rect 18679 -1522 18695 -1470
rect 18747 -1522 18763 -1470
rect 18815 -1522 18831 -1470
rect 18883 -1522 18899 -1470
rect 18951 -1522 18967 -1470
rect 19019 -1522 19035 -1470
rect 19087 -1522 19103 -1470
rect 19155 -1522 19171 -1470
rect 19223 -1522 19229 -1470
rect 20190 -1522 20196 -1470
rect 20248 -1522 20264 -1470
rect 20316 -1522 20332 -1470
rect 20384 -1522 20400 -1470
rect 20452 -1522 20468 -1470
rect 20520 -1522 20536 -1470
rect 20588 -1522 20604 -1470
rect 20656 -1522 20672 -1470
rect 20724 -1522 20740 -1470
rect 20792 -1522 20808 -1470
rect 20860 -1522 20876 -1470
rect 20928 -1522 20944 -1470
rect 20996 -1522 21012 -1470
rect 21064 -1522 21070 -1470
tri 13632 -1604 13714 -1522 se
rect 13714 -1604 14594 -1522
tri 14594 -1604 14676 -1522 sw
tri 18267 -1604 18349 -1522 se
rect 18349 -1604 19229 -1522
tri 19229 -1604 19311 -1522 sw
tri 20108 -1604 20190 -1522 se
rect 20190 -1604 21070 -1522
tri 21070 -1604 21152 -1522 sw
tri 13628 -1608 13632 -1604 se
rect 13632 -1608 14676 -1604
tri 14676 -1608 14680 -1604 sw
tri 18263 -1608 18267 -1604 se
rect 18267 -1608 19311 -1604
tri 19311 -1608 19315 -1604 sw
tri 20104 -1608 20108 -1604 se
rect 20108 -1608 21152 -1604
tri 21152 -1608 21156 -1604 sw
tri 26695 -1608 26699 -1604 se
rect 26699 -1608 26827 -1604
tri 26827 -1608 26831 -1604 sw
rect 684 -1792 930 -1613
rect 26238 -1798 26443 -1608
rect 26695 -1798 26831 -1608
tri 26238 -1802 26242 -1798 ne
rect 26242 -1802 26439 -1798
tri 26439 -1802 26443 -1798 nw
rect 1309 -6932 6121 -6931
tri 6121 -6932 6122 -6931 sw
rect 1309 -6934 6142 -6932
tri 6142 -6934 6144 -6932 sw
tri 2956 -7172 2958 -7170 ne
rect 2958 -7172 3011 -6934
tri 12399 -6941 12400 -6940 se
rect 12400 -6941 12401 -6940
tri 6650 -6944 6653 -6941 se
rect 6653 -6944 6700 -6941
tri 12396 -6944 12399 -6941 se
rect 12399 -6944 12401 -6941
tri 6642 -6952 6650 -6944 se
rect 6650 -6952 6700 -6944
rect 6421 -7142 6700 -6952
tri 6596 -7143 6597 -7142 ne
rect 6597 -7143 6700 -7142
rect 6756 -7075 6762 -7023
rect 6814 -7075 6829 -7023
rect 6881 -7075 6896 -7023
rect 6948 -7075 6963 -7023
rect 7015 -7075 7030 -7023
rect 7082 -7075 7096 -7023
rect 7148 -7075 7154 -7023
rect 6756 -7091 7154 -7075
rect 6756 -7143 6762 -7091
rect 6814 -7143 6829 -7091
rect 6881 -7143 6896 -7091
rect 6948 -7143 6963 -7091
rect 7015 -7143 7030 -7091
rect 7082 -7143 7096 -7091
rect 7148 -7143 7154 -7091
tri 6152 -7204 6184 -7172 ne
tri 6236 -7204 6268 -7172 nw
rect 12308 -7217 12311 -7211
tri 12311 -7217 12317 -7211 nw
rect 10222 -7230 10257 -7217
tri 10257 -7230 10270 -7217 nw
tri 6318 -7255 6343 -7230 ne
rect 6343 -7255 6395 -7230
tri 6395 -7239 6404 -7230 nw
rect 10222 -7239 10248 -7230
tri 10248 -7239 10257 -7230 nw
rect 10222 -7255 10232 -7239
tri 10232 -7255 10248 -7239 nw
tri 10222 -7265 10232 -7255 nw
rect 8484 -7288 8507 -7273
tri 8507 -7288 8522 -7273 nw
tri 9101 -7288 9116 -7273 ne
rect 9116 -7288 9125 -7273
tri 6012 -7293 6017 -7288 se
rect 6017 -7293 6047 -7288
rect 6012 -7339 6047 -7293
rect 8484 -7297 8498 -7288
tri 8498 -7297 8507 -7288 nw
tri 9116 -7297 9125 -7288 ne
rect 8484 -7299 8496 -7297
tri 8496 -7299 8498 -7297 nw
tri 7090 -7307 7098 -7299 ne
rect 7098 -7307 7116 -7299
rect 8484 -7305 8490 -7299
tri 8490 -7305 8496 -7299 nw
tri 10334 -7305 10340 -7299 se
rect 8484 -7310 8485 -7305
tri 8485 -7310 8490 -7305 nw
tri 10329 -7310 10334 -7305 se
rect 10334 -7310 10340 -7305
tri 10320 -7319 10329 -7310 se
rect 10329 -7319 10340 -7310
tri 6012 -7340 6013 -7339 ne
rect 6013 -7340 6047 -7339
rect 9922 -7328 9924 -7319
tri 9924 -7328 9933 -7319 sw
tri 10311 -7328 10320 -7319 se
rect 10320 -7328 10340 -7319
rect 11142 -7328 11149 -7305
tri 11149 -7328 11172 -7305 nw
tri 1414 -7365 1434 -7345 se
tri 1897 -7351 1903 -7345 se
rect 1903 -7351 1949 -7345
tri 1643 -7364 1656 -7351 se
tri 1387 -7392 1414 -7365 se
rect 1414 -7392 1434 -7365
tri 1385 -7394 1387 -7392 se
rect 1387 -7394 1434 -7392
tri 1480 -7365 1481 -7364 sw
tri 1642 -7365 1643 -7364 se
rect 1643 -7365 1656 -7364
rect 1480 -7392 1481 -7365
tri 1481 -7392 1508 -7365 sw
tri 1619 -7388 1642 -7365 se
rect 1642 -7388 1656 -7365
rect 1897 -7353 1949 -7351
tri 1949 -7353 1957 -7345 sw
rect 1897 -7388 1977 -7353
rect 9922 -7359 9933 -7328
tri 11142 -7335 11149 -7328 nw
rect 9922 -7363 9929 -7359
tri 9929 -7363 9933 -7359 nw
tri 10336 -7363 10340 -7359 ne
rect 10340 -7363 10341 -7359
rect 9922 -7365 9927 -7363
tri 9927 -7365 9929 -7363 nw
tri 1615 -7392 1619 -7388 se
rect 1619 -7392 1656 -7388
rect 1480 -7394 1508 -7392
tri 1508 -7394 1510 -7392 sw
tri 1613 -7394 1615 -7392 se
rect 1615 -7394 1656 -7392
rect 1860 -7397 1977 -7388
tri 3260 -7392 3284 -7368 se
rect 3284 -7392 3304 -7368
tri 3258 -7394 3260 -7392 se
rect 3260 -7394 3304 -7392
tri 12162 -7394 12164 -7392 se
tri 12164 -7394 12166 -7392 sw
rect 3150 -7396 3304 -7394
tri 1977 -7397 1978 -7396 nw
rect 1702 -7401 1741 -7397
tri 1741 -7401 1745 -7397 nw
tri 1860 -7401 1864 -7397 ne
rect 1864 -7401 1903 -7397
rect 1702 -7426 1716 -7401
tri 1716 -7426 1741 -7401 nw
tri 1864 -7426 1889 -7401 ne
rect 1889 -7426 1903 -7401
rect 1949 -7401 1973 -7397
tri 1973 -7401 1977 -7397 nw
tri 1949 -7425 1973 -7401 nw
tri 1702 -7440 1716 -7426 nw
tri 1889 -7440 1903 -7426 ne
rect 3150 -7440 3164 -7396
tri 1399 -7445 1404 -7440 ne
rect 1404 -7445 1434 -7440
tri 1404 -7456 1415 -7445 ne
rect 1415 -7456 1434 -7445
tri 1415 -7475 1434 -7456 ne
rect 1480 -7445 1510 -7440
tri 1510 -7445 1515 -7440 nw
tri 3150 -7445 3155 -7440 ne
rect 3155 -7445 3164 -7440
rect 1480 -7456 1499 -7445
tri 1499 -7456 1510 -7445 nw
tri 3155 -7448 3158 -7445 ne
rect 3158 -7448 3164 -7445
rect 3216 -7448 3228 -7396
rect 3280 -7448 3304 -7396
tri 7663 -7426 7688 -7401 se
rect 7688 -7426 7694 -7401
tri 3243 -7456 3251 -7448 ne
rect 3251 -7456 3304 -7448
tri 9295 -7456 9306 -7445 se
tri 1480 -7475 1499 -7456 nw
tri 3251 -7475 3270 -7456 ne
rect 3270 -7475 3304 -7456
tri 3270 -7481 3276 -7475 ne
rect 3276 -7481 3304 -7475
tri 7849 -7481 7874 -7456 se
rect 7874 -7481 7880 -7456
tri 9270 -7481 9295 -7456 se
rect 9295 -7481 9306 -7456
rect 12641 -7453 12647 -7401
rect 12699 -7453 12739 -7401
rect 12791 -7453 12831 -7401
rect 12883 -7453 12922 -7401
rect 12974 -7453 13013 -7401
rect 13065 -7453 13071 -7401
tri 3276 -7489 3284 -7481 ne
rect 3284 -7489 3304 -7481
tri 1967 -7509 1984 -7492 se
rect 12641 -7505 13071 -7453
tri 1943 -7533 1967 -7509 se
rect 1967 -7533 1984 -7509
tri 6160 -7533 6184 -7509 se
tri 6157 -7536 6160 -7533 se
rect 6160 -7536 6184 -7533
rect 121 -7564 122 -7537
tri 122 -7564 149 -7537 nw
rect 12641 -7557 12647 -7505
rect 12699 -7557 12739 -7505
rect 12791 -7557 12831 -7505
rect 12883 -7557 12922 -7505
rect 12974 -7557 13013 -7505
rect 13065 -7557 13071 -7505
tri 121 -7565 122 -7564 nw
tri 3103 -7565 3104 -7564 se
rect 3104 -7565 3142 -7564
tri 3102 -7566 3103 -7565 se
rect 3103 -7566 3142 -7565
tri 1975 -7575 1984 -7566 ne
rect 1984 -7575 1987 -7566
tri 3093 -7575 3102 -7566 se
rect 3102 -7575 3142 -7566
tri 3080 -7588 3093 -7575 se
rect 3093 -7588 3142 -7575
tri 3071 -7597 3080 -7588 se
rect 3080 -7597 3142 -7588
tri 6159 -7597 6168 -7588 ne
rect 6168 -7597 6184 -7588
tri 3057 -7611 3071 -7597 se
rect 3071 -7611 3142 -7597
rect 3057 -7613 3142 -7611
tri 3142 -7613 3158 -7597 sw
tri 6168 -7613 6184 -7597 ne
rect 12641 -7609 13071 -7557
rect 3057 -7622 3158 -7613
tri 3158 -7622 3167 -7613 sw
rect 3057 -7633 3167 -7622
tri 3057 -7649 3073 -7633 ne
rect 3073 -7649 3167 -7633
tri 1863 -7680 1894 -7649 ne
rect 1894 -7655 1948 -7649
tri 1948 -7655 1954 -7649 nw
tri 3073 -7655 3079 -7649 ne
rect 3079 -7655 3167 -7649
rect 1894 -7661 1942 -7655
tri 1942 -7661 1948 -7655 nw
tri 3079 -7661 3085 -7655 ne
rect 3085 -7661 3167 -7655
tri 6178 -7661 6184 -7655 se
rect 1894 -7672 1931 -7661
tri 1931 -7672 1942 -7661 nw
tri 3085 -7672 3096 -7661 ne
rect 1894 -7677 1926 -7672
tri 1926 -7677 1931 -7672 nw
rect 3096 -7674 3167 -7661
tri 6165 -7674 6178 -7661 se
rect 6178 -7674 6184 -7661
rect 8279 -7667 8285 -7615
rect 8337 -7667 8377 -7615
rect 8429 -7667 8469 -7615
rect 8521 -7667 8527 -7615
rect 12641 -7661 12647 -7609
rect 12699 -7661 12739 -7609
rect 12791 -7661 12831 -7609
rect 12883 -7661 12922 -7609
rect 12974 -7661 13013 -7609
rect 13065 -7661 13071 -7609
rect 3096 -7677 3142 -7674
tri 3142 -7677 3145 -7674 nw
tri 6162 -7677 6165 -7674 se
rect 6165 -7677 6184 -7674
rect 1894 -7680 1923 -7677
tri 1923 -7680 1926 -7677 nw
tri 6159 -7680 6162 -7677 se
rect 6162 -7680 6184 -7677
tri 5617 -7683 5620 -7680 se
rect 5620 -7683 5714 -7680
tri 621 -7684 622 -7683 se
rect 622 -7684 627 -7683
tri 1642 -7684 1643 -7683 se
rect 1643 -7684 1771 -7683
tri 618 -7687 621 -7684 se
rect 621 -7687 627 -7684
rect 618 -7733 627 -7687
tri 618 -7735 620 -7733 ne
rect 620 -7735 627 -7733
tri 883 -7687 886 -7684 se
rect 883 -7733 886 -7687
tri 883 -7735 885 -7733 ne
rect 885 -7735 886 -7733
tri 885 -7736 886 -7735 ne
tri 1158 -7686 1160 -7684 sw
tri 1640 -7686 1642 -7684 se
rect 1642 -7686 1771 -7684
tri 1771 -7686 1774 -7683 sw
tri 5614 -7686 5617 -7683 se
rect 5617 -7686 5714 -7683
tri 6153 -7686 6159 -7680 se
rect 6159 -7686 6184 -7680
rect 1158 -7687 1160 -7686
tri 1160 -7687 1161 -7686 sw
rect 1158 -7733 1161 -7687
rect 1158 -7735 1159 -7733
tri 1159 -7735 1161 -7733 nw
tri 1639 -7687 1640 -7686 se
rect 1640 -7687 1774 -7686
tri 1774 -7687 1775 -7686 sw
rect 1639 -7731 1775 -7687
tri 5613 -7687 5614 -7686 se
rect 5614 -7687 5714 -7686
tri 2639 -7721 2651 -7709 se
rect 2651 -7721 2779 -7709
tri 2779 -7721 2791 -7709 sw
rect 1639 -7733 1773 -7731
tri 1773 -7733 1775 -7731 nw
tri 2638 -7722 2639 -7721 se
rect 2639 -7722 2791 -7721
tri 2791 -7722 2792 -7721 sw
tri 1639 -7735 1641 -7733 ne
rect 1641 -7735 1771 -7733
tri 1771 -7735 1773 -7733 nw
tri 1158 -7736 1159 -7735 nw
rect 2638 -7761 2792 -7722
tri 3214 -7724 3217 -7721 se
rect 3217 -7724 3219 -7721
rect 3214 -7766 3219 -7724
rect 5613 -7731 5714 -7687
rect 5613 -7733 5712 -7731
tri 5712 -7733 5714 -7731 nw
rect 8946 -7762 8948 -7737
tri 8948 -7762 8973 -7737 nw
tri 9683 -7762 9708 -7737 ne
tri 8946 -7764 8948 -7762 nw
rect 3214 -7768 3217 -7766
tri 3217 -7768 3219 -7766 nw
tri 4173 -7768 4175 -7766 ne
rect 4175 -7768 4403 -7766
tri 6574 -7808 6609 -7773 sw
tri 8362 -7832 8374 -7820 ne
rect 8374 -7832 8397 -7820
tri 3442 -7864 3474 -7832 ne
rect 3474 -7864 3479 -7832
tri 8374 -7851 8393 -7832 ne
rect 8393 -7851 8397 -7832
rect 8449 -7830 8470 -7820
tri 8470 -7830 8480 -7820 nw
rect 8449 -7832 8468 -7830
tri 8468 -7832 8470 -7830 nw
tri 9667 -7832 9669 -7830 sw
tri 10806 -7832 10808 -7830 se
tri 8449 -7851 8468 -7832 nw
tri 8393 -7855 8397 -7851 ne
rect 9667 -7855 9669 -7832
tri 9669 -7855 9692 -7832 sw
tri 10783 -7855 10806 -7832 se
rect 10806 -7855 10808 -7832
tri 3474 -7869 3479 -7864 ne
tri 8226 -7869 8231 -7864 ne
rect 8231 -7869 8260 -7864
tri 8231 -7898 8260 -7869 ne
tri 8390 -7898 8397 -7891 se
tri 8388 -7900 8390 -7898 se
rect 8390 -7900 8397 -7898
tri 9402 -7900 9404 -7898 sw
tri 8367 -7921 8388 -7900 se
rect 8388 -7921 8397 -7900
tri 8449 -7921 8470 -7900 sw
rect 9402 -7921 9404 -7900
tri 9404 -7921 9425 -7900 sw
rect 9402 -7923 9425 -7921
tri 9425 -7923 9427 -7921 sw
rect 5467 -7973 5545 -7966
tri 5545 -7973 5552 -7966 sw
rect 5467 -7978 5552 -7973
tri 5552 -7978 5557 -7973 sw
tri 8602 -7978 8607 -7973 se
tri 5463 -7984 5467 -7980 se
rect 5467 -7984 5557 -7978
tri 1386 -8019 1421 -7984 nw
tri 5449 -7998 5463 -7984 se
rect 5463 -7997 5557 -7984
tri 5557 -7997 5576 -7978 sw
tri 8583 -7997 8602 -7978 se
rect 8602 -7997 8607 -7978
tri 9253 -7997 9272 -7978 sw
rect 5463 -7998 5576 -7997
rect 5449 -8002 5576 -7998
tri 5576 -8002 5581 -7997 sw
tri 8578 -8002 8583 -7997 se
rect 8583 -8002 8607 -7997
tri 2028 -8068 2067 -8029 se
rect 2067 -8068 2072 -8029
rect 5449 -8044 5581 -8002
tri 5581 -8044 5623 -8002 sw
rect 5449 -8048 5623 -8044
tri 5623 -8048 5627 -8044 sw
tri 8256 -8048 8260 -8044 se
rect 5449 -8050 5601 -8048
tri 5449 -8061 5460 -8050 ne
rect 5460 -8061 5601 -8050
tri 2012 -8084 2028 -8068 se
rect 2028 -8084 2072 -8068
rect 2136 -8068 2158 -8061
tri 2158 -8068 2165 -8061 nw
tri 5460 -8068 5467 -8061 ne
rect 5467 -8068 5601 -8061
rect 2136 -8084 2142 -8068
tri 2142 -8084 2158 -8068 nw
tri 2136 -8090 2142 -8084 nw
rect 5519 -8100 5601 -8068
tri 8226 -8078 8256 -8048 se
rect 8256 -8078 8260 -8048
tri 11993 -8078 12004 -8067 ne
rect 12004 -8078 12021 -8067
tri 12004 -8092 12018 -8078 ne
rect 12018 -8092 12021 -8078
rect 5519 -8114 5537 -8100
tri 5537 -8114 5551 -8100 nw
rect 10695 -8114 10784 -8092
tri 12018 -8095 12021 -8092 ne
rect 12067 -8078 12084 -8067
tri 12084 -8078 12095 -8067 nw
tri 12067 -8095 12084 -8078 nw
rect 5519 -8121 5530 -8114
tri 5530 -8121 5537 -8114 nw
tri 10675 -8121 10682 -8114 se
rect 10682 -8121 10800 -8114
tri 10800 -8121 10803 -8118 sw
tri 5519 -8132 5530 -8121 nw
tri 2944 -8145 2952 -8137 ne
rect 2952 -8145 3080 -8137
tri 3080 -8145 3088 -8137 nw
rect 10423 -8162 10487 -8124
rect 10695 -8146 10784 -8121
tri 6255 -8194 6271 -8178 ne
rect 6271 -8194 6285 -8178
tri 9530 -8183 9533 -8180 sw
tri 1386 -8206 1398 -8194 sw
tri 1681 -8206 1693 -8194 se
tri 1317 -8229 1340 -8206 se
rect 1386 -8229 1398 -8206
tri 1398 -8229 1421 -8206 sw
tri 1658 -8229 1681 -8206 se
rect 1681 -8229 1693 -8206
tri 1739 -8203 1748 -8194 sw
tri 6271 -8203 6280 -8194 ne
rect 6280 -8203 6285 -8194
rect 1739 -8208 1748 -8203
tri 1748 -8208 1753 -8203 sw
tri 5110 -8208 5115 -8203 ne
rect 5115 -8208 5135 -8203
tri 6280 -8208 6285 -8203 ne
tri 8636 -8187 8640 -8183 sw
rect 9530 -8187 9533 -8183
tri 9533 -8187 9537 -8183 sw
rect 8636 -8194 8640 -8187
tri 8640 -8194 8647 -8187 sw
tri 8899 -8194 8906 -8187 se
rect 9530 -8194 9537 -8187
tri 9537 -8194 9544 -8187 sw
rect 8636 -8208 8647 -8194
tri 8647 -8208 8661 -8194 sw
tri 8885 -8208 8899 -8194 se
rect 8899 -8208 8906 -8194
rect 1739 -8226 1753 -8208
tri 1753 -8226 1771 -8208 sw
tri 5115 -8226 5133 -8208 ne
rect 5133 -8226 5135 -8208
rect 8636 -8214 8661 -8208
tri 8661 -8214 8667 -8208 sw
tri 8879 -8214 8885 -8208 se
rect 8885 -8214 8906 -8208
rect 1739 -8228 1771 -8226
tri 1771 -8228 1773 -8226 sw
tri 5133 -8228 5135 -8226 ne
tri 8226 -8228 8228 -8226 ne
rect 8228 -8228 8260 -8226
rect 1739 -8229 1773 -8228
tri 1773 -8229 1774 -8228 sw
tri 8228 -8229 8229 -8228 ne
rect 8229 -8229 8260 -8228
tri 8229 -8238 8238 -8229 ne
rect 8238 -8238 8260 -8229
tri 5863 -8260 5885 -8238 sw
tri 8238 -8260 8260 -8238 ne
rect 8636 -8254 8667 -8214
rect 11829 -8226 11889 -8194
tri 12407 -8226 12408 -8225 sw
tri 10836 -8227 10837 -8226 ne
rect 10837 -8227 10980 -8226
tri 9064 -8252 9089 -8227 sw
tri 10837 -8252 10862 -8227 ne
rect 10862 -8252 10980 -8227
tri 10980 -8252 11006 -8226 nw
rect 9064 -8253 9089 -8252
tri 9089 -8253 9090 -8252 sw
rect 12407 -8253 12408 -8226
tri 12408 -8253 12435 -8226 sw
rect 9064 -8254 9090 -8253
tri 9090 -8254 9091 -8253 sw
rect 8636 -8260 8661 -8254
tri 8661 -8260 8667 -8254 nw
rect 5863 -8284 5885 -8260
tri 5885 -8284 5909 -8260 sw
rect 8636 -8284 8637 -8260
tri 8637 -8284 8661 -8260 nw
tri 4525 -8308 4549 -8284 ne
rect 4549 -8308 4699 -8284
tri 4699 -8308 4723 -8284 nw
rect 5863 -8285 5909 -8284
tri 5909 -8285 5910 -8284 sw
tri 8636 -8285 8637 -8284 nw
tri 4549 -8318 4559 -8308 ne
rect 4559 -8318 4689 -8308
tri 4689 -8318 4699 -8308 nw
rect 5145 -8337 5151 -8285
rect 5203 -8337 5250 -8285
rect 5302 -8337 5348 -8285
rect 5400 -8337 5406 -8285
rect 5863 -8286 5910 -8285
tri 5910 -8286 5911 -8285 sw
rect 5863 -8287 5911 -8286
tri 5911 -8287 5912 -8286 sw
tri 1974 -8360 1989 -8345 ne
rect 1989 -8360 2008 -8345
tri 1989 -8373 2002 -8360 ne
rect 2002 -8373 2008 -8360
tri 2002 -8376 2005 -8373 ne
rect 2005 -8376 2008 -8373
rect 5145 -8359 5406 -8337
rect 5145 -8411 5151 -8359
rect 5203 -8411 5250 -8359
rect 5302 -8411 5348 -8359
rect 5400 -8411 5406 -8359
rect 5145 -8433 5406 -8411
rect 5145 -8485 5151 -8433
rect 5203 -8485 5250 -8433
rect 5302 -8485 5348 -8433
rect 5400 -8485 5406 -8433
rect 5591 -8339 5597 -8287
rect 5649 -8339 5662 -8287
rect 5591 -8351 5662 -8339
rect 5591 -8403 5597 -8351
rect 5649 -8403 5662 -8351
rect 5591 -8415 5662 -8403
rect 5591 -8467 5597 -8415
rect 5649 -8467 5662 -8415
rect 5906 -8467 5912 -8287
tri 9882 -8300 9896 -8286 ne
tri 8034 -8311 8037 -8308 se
rect 8037 -8311 8131 -8308
rect 7639 -8357 7738 -8311
rect 8034 -8357 8131 -8311
tri 8034 -8360 8037 -8357 ne
rect 8037 -8360 8131 -8357
rect 8737 -8406 8738 -8373
tri 8738 -8406 8771 -8373 nw
tri 8259 -8407 8260 -8406 se
tri 8737 -8407 8738 -8406 nw
tri 8226 -8440 8259 -8407 se
rect 8259 -8440 8260 -8407
rect 5863 -8496 5883 -8467
tri 5883 -8496 5912 -8467 nw
rect 8845 -8457 8915 -8454
tri 8915 -8457 8918 -8454 sw
tri 5457 -8506 5467 -8496 se
tri 5453 -8510 5457 -8506 se
rect 5457 -8510 5467 -8506
tri 5427 -8536 5453 -8510 se
rect 5453 -8536 5467 -8510
rect 5863 -8506 5873 -8496
tri 5873 -8506 5883 -8496 nw
rect 8845 -8503 8918 -8457
rect 8845 -8506 8915 -8503
tri 8915 -8506 8918 -8503 nw
rect 5863 -8510 5869 -8506
tri 5869 -8510 5873 -8506 nw
tri 5863 -8516 5869 -8510 nw
tri 6218 -8516 6224 -8510 se
tri 6198 -8536 6218 -8516 se
rect 6218 -8536 6224 -8516
tri 6190 -8544 6198 -8536 se
rect 6198 -8544 6224 -8536
tri 8737 -8569 8753 -8553 sw
tri 5588 -8572 5591 -8569 se
rect 5591 -8572 5647 -8569
tri 1128 -8578 1134 -8572 sw
tri 5582 -8578 5588 -8572 se
rect 5588 -8578 5647 -8572
tri 964 -8612 998 -8578 se
rect 1128 -8581 1134 -8578
tri 1134 -8581 1137 -8578 sw
tri 5579 -8581 5582 -8578 se
rect 5582 -8581 5647 -8578
rect 1128 -8582 1137 -8581
tri 1137 -8582 1138 -8581 sw
tri 1923 -8582 1924 -8581 ne
rect 1924 -8582 2132 -8581
tri 5578 -8582 5579 -8581 se
rect 5579 -8582 5647 -8581
rect 1128 -8587 1138 -8582
tri 1138 -8587 1143 -8582 sw
tri 5573 -8587 5578 -8582 se
rect 5578 -8587 5647 -8582
rect 8737 -8587 8753 -8569
tri 8753 -8587 8771 -8569 sw
rect 1128 -8592 1143 -8587
tri 1143 -8592 1148 -8587 sw
tri 5568 -8592 5573 -8587 se
rect 5573 -8592 5647 -8587
rect 1128 -8593 1148 -8592
tri 1148 -8593 1149 -8592 sw
tri 5567 -8593 5568 -8592 se
rect 5568 -8593 5647 -8592
tri 6318 -8593 6319 -8592 se
rect 1128 -8612 1149 -8593
tri 1149 -8612 1168 -8593 sw
tri 5548 -8612 5567 -8593 se
rect 5567 -8612 5647 -8593
tri 5545 -8615 5548 -8612 se
rect 5548 -8615 5647 -8612
tri 6296 -8615 6318 -8593 se
rect 6318 -8615 6319 -8593
tri 6287 -8624 6296 -8615 se
rect 6296 -8624 6319 -8615
tri 6371 -8624 6402 -8593 sw
tri 11969 -8679 12003 -8645 ne
rect 8527 -8688 8546 -8687
tri 8546 -8688 8547 -8687 sw
tri 8468 -8720 8500 -8688 se
rect 8500 -8720 8547 -8688
tri 8547 -8720 8579 -8688 sw
tri 11965 -8801 12003 -8763 se
tri 13207 -8842 13241 -8808 se
rect 6756 -8917 6762 -8865
rect 6814 -8917 6829 -8865
rect 6881 -8917 6896 -8865
rect 6948 -8917 6963 -8865
rect 7015 -8917 7030 -8865
rect 7082 -8917 7096 -8865
rect 7148 -8917 7154 -8865
rect 6756 -8933 7154 -8917
rect 6756 -8960 6762 -8933
tri 6731 -8984 6755 -8960 ne
rect 6755 -8984 6762 -8960
tri 6755 -8985 6756 -8984 ne
rect 6756 -8985 6762 -8984
rect 6814 -8985 6829 -8933
rect 6881 -8985 6896 -8933
rect 6948 -8985 6963 -8933
rect 7015 -8985 7030 -8933
rect 7082 -8985 7096 -8933
rect 7148 -8960 7154 -8933
rect 9440 -8960 9464 -8959
tri 9464 -8960 9465 -8959 nw
rect 7148 -8984 7155 -8960
tri 7155 -8984 7179 -8960 nw
tri 8735 -8984 8759 -8960 ne
tri 9440 -8984 9464 -8960 nw
rect 7148 -8985 7154 -8984
tri 7154 -8985 7155 -8984 nw
<< rmetal1 >>
rect 23654 2858 23734 2860
rect 23811 2731 23813 2811
<< via1 >>
rect 804 15831 856 15883
rect 888 15831 940 15883
rect 972 15831 1024 15883
rect 804 15752 856 15804
rect 888 15752 940 15804
rect 972 15752 1024 15804
rect 804 15673 856 15725
rect 888 15673 940 15725
rect 972 15673 1024 15725
rect 804 15594 856 15646
rect 888 15594 940 15646
rect 972 15594 1024 15646
rect 25109 7348 25225 7353
rect 23031 7320 23083 7329
rect 23031 7286 23037 7320
rect 23037 7286 23071 7320
rect 23071 7286 23083 7320
rect 23031 7277 23083 7286
rect 23097 7320 23149 7329
rect 23097 7286 23109 7320
rect 23109 7286 23143 7320
rect 23143 7286 23149 7320
rect 23097 7277 23149 7286
rect 25109 7242 25115 7348
rect 25115 7242 25221 7348
rect 25221 7242 25225 7348
rect 25109 7237 25225 7242
rect 23013 7117 23065 7122
rect 23013 7083 23019 7117
rect 23019 7083 23053 7117
rect 23053 7083 23065 7117
rect 23013 7070 23065 7083
rect 23013 7045 23065 7058
rect 23013 7011 23019 7045
rect 23019 7011 23053 7045
rect 23053 7011 23065 7045
rect 23013 7006 23065 7011
rect 25105 7116 25221 7122
rect 25105 7010 25106 7116
rect 25106 7010 25212 7116
rect 25212 7010 25221 7116
rect 25105 7006 25221 7010
rect 6339 6480 6391 6532
rect 6405 6480 6457 6532
rect 6471 6480 6523 6532
rect 6537 6480 6589 6532
rect 6603 6480 6655 6532
rect 6668 6480 6720 6532
rect 6733 6480 6785 6532
rect 6798 6480 6850 6532
rect 6863 6480 6915 6532
rect 6928 6480 6980 6532
rect 6993 6480 7045 6532
rect 7058 6480 7110 6532
rect 7123 6480 7175 6532
rect 7188 6480 7240 6532
rect 7253 6480 7305 6532
rect 7318 6480 7370 6532
rect 7383 6480 7435 6532
rect 7448 6480 7500 6532
rect 7513 6480 7565 6532
rect 7578 6480 7630 6532
rect 6339 6364 6391 6416
rect 6405 6364 6457 6416
rect 6471 6364 6523 6416
rect 6537 6364 6589 6416
rect 6603 6364 6655 6416
rect 6668 6364 6720 6416
rect 6733 6364 6785 6416
rect 6798 6364 6850 6416
rect 6863 6364 6915 6416
rect 6928 6364 6980 6416
rect 6993 6364 7045 6416
rect 7058 6364 7110 6416
rect 7123 6364 7175 6416
rect 7188 6364 7240 6416
rect 7253 6364 7305 6416
rect 7318 6364 7370 6416
rect 7383 6364 7435 6416
rect 7448 6364 7500 6416
rect 7513 6364 7565 6416
rect 7578 6364 7630 6416
rect 18359 6480 18411 6532
rect 18428 6480 18480 6532
rect 18497 6480 18549 6532
rect 18565 6480 18617 6532
rect 18633 6480 18685 6532
rect 18701 6480 18753 6532
rect 18769 6480 18821 6532
rect 18837 6480 18889 6532
rect 18905 6480 18957 6532
rect 18973 6480 19025 6532
rect 19041 6480 19093 6532
rect 19109 6480 19161 6532
rect 19177 6480 19229 6532
rect 18359 6364 18411 6416
rect 18428 6364 18480 6416
rect 18497 6364 18549 6416
rect 18565 6364 18617 6416
rect 18633 6364 18685 6416
rect 18701 6364 18753 6416
rect 18769 6364 18821 6416
rect 18837 6364 18889 6416
rect 18905 6364 18957 6416
rect 18973 6364 19025 6416
rect 19041 6364 19093 6416
rect 19109 6364 19161 6416
rect 19177 6364 19229 6416
rect 20198 6480 20250 6532
rect 20267 6480 20319 6532
rect 20336 6480 20388 6532
rect 20404 6480 20456 6532
rect 20472 6480 20524 6532
rect 20540 6480 20592 6532
rect 20608 6480 20660 6532
rect 20676 6480 20728 6532
rect 20744 6480 20796 6532
rect 20812 6480 20864 6532
rect 20880 6480 20932 6532
rect 20948 6480 21000 6532
rect 21016 6480 21068 6532
rect 20198 6364 20250 6416
rect 20267 6364 20319 6416
rect 20336 6364 20388 6416
rect 20404 6364 20456 6416
rect 20472 6364 20524 6416
rect 20540 6364 20592 6416
rect 20608 6364 20660 6416
rect 20676 6364 20728 6416
rect 20744 6364 20796 6416
rect 20812 6364 20864 6416
rect 20880 6364 20932 6416
rect 20948 6364 21000 6416
rect 21016 6364 21068 6416
rect 22981 6480 23033 6532
rect 23072 6480 23124 6532
rect 22981 6364 23033 6416
rect 23072 6364 23124 6416
rect 23154 5593 23270 5773
rect 8094 5498 8146 5550
rect 8158 5498 8210 5550
rect 11314 5498 11366 5550
rect 11378 5498 11430 5550
rect 14534 5498 14586 5550
rect 14598 5498 14650 5550
rect 17754 5498 17806 5550
rect 17818 5498 17870 5550
rect 20974 5498 21026 5550
rect 21038 5498 21090 5550
rect 24194 5498 24246 5550
rect 24258 5498 24310 5550
rect 6127 5387 6179 5439
rect 6191 5387 6243 5439
rect 3041 5312 3093 5364
rect 3105 5312 3157 5364
rect 25583 5323 25699 5439
rect 2441 5190 2493 5242
rect 2505 5190 2557 5242
rect 16270 5165 16322 5217
rect 16337 5165 16389 5217
rect 16404 5165 16456 5217
rect 16470 5165 16522 5217
rect 23353 5166 23469 5282
rect 24798 5214 24850 5266
rect 24862 5214 24914 5266
rect 25842 5166 25958 5282
rect 2514 5103 2566 5155
rect 2578 5103 2630 5155
rect 6280 4966 6332 5018
rect 6344 4966 6396 5018
rect 7638 4966 7690 5018
rect 7702 4966 7754 5018
rect 5429 4888 5481 4940
rect 5507 4888 5559 4940
rect 5585 4888 5637 4940
rect 7839 4888 7891 4940
rect 7908 4888 7960 4940
rect 7976 4888 8028 4940
rect 13450 4888 13502 4940
rect 13519 4888 13571 4940
rect 13587 4888 13639 4940
rect 16270 4888 16322 4940
rect 16337 4888 16389 4940
rect 16404 4888 16456 4940
rect 16470 4888 16522 4940
rect 19519 4888 19571 4940
rect 19588 4888 19640 4940
rect 19656 4888 19708 4940
rect 22913 4888 22965 4940
rect 22982 4888 23034 4940
rect 23050 4888 23102 4940
rect 2686 4734 2738 4786
rect 2750 4734 2802 4786
rect 22913 4574 22965 4626
rect 22982 4574 23034 4626
rect 23050 4574 23102 4626
rect 19519 4514 19571 4566
rect 19588 4514 19640 4566
rect 19656 4514 19708 4566
rect 7839 4454 7891 4506
rect 7908 4454 7960 4506
rect 7976 4454 8028 4506
rect 8092 4454 8144 4506
rect 8156 4454 8208 4506
rect 8698 4454 8750 4506
rect 8762 4454 8814 4506
rect 11918 4454 11970 4506
rect 11982 4454 12034 4506
rect 13219 4454 13271 4506
rect 13283 4454 13335 4506
rect 13787 4454 13839 4506
rect 13851 4454 13903 4506
rect 15138 4454 15190 4506
rect 15202 4454 15254 4506
rect 18358 4454 18410 4506
rect 18422 4454 18474 4506
rect 19299 4454 19351 4506
rect 19363 4454 19415 4506
rect 19867 4454 19919 4506
rect 19931 4454 19983 4506
rect 21578 4454 21630 4506
rect 21642 4454 21694 4506
rect 22636 4454 22688 4506
rect 22700 4454 22752 4506
rect 23663 4500 23779 4616
rect 25742 4544 25858 4660
rect 13450 4392 13502 4444
rect 13519 4392 13571 4444
rect 13587 4392 13639 4444
rect 2844 2418 2896 2470
rect 2995 2418 3047 2470
rect 2844 2354 2896 2406
rect 2995 2354 3047 2406
rect 2326 1706 2378 1758
rect 2844 1706 2896 1758
rect 2326 1642 2378 1694
rect 2844 1642 2896 1694
rect 23720 1228 23772 1280
rect 23720 1164 23772 1216
rect 23720 1100 23772 1152
rect 2850 696 2902 748
rect 2914 696 2966 748
rect 2850 -72 2902 -20
rect 2914 -72 2966 -20
rect 2163 -533 2215 -481
rect 2227 -533 2279 -481
rect 23674 -533 23726 -481
rect 23738 -533 23790 -481
rect 23802 -533 23854 -481
rect 13720 -1522 13772 -1470
rect 13788 -1522 13840 -1470
rect 13856 -1522 13908 -1470
rect 13924 -1522 13976 -1470
rect 13992 -1522 14044 -1470
rect 14060 -1522 14112 -1470
rect 14128 -1522 14180 -1470
rect 14196 -1522 14248 -1470
rect 14264 -1522 14316 -1470
rect 14332 -1522 14384 -1470
rect 14400 -1522 14452 -1470
rect 14468 -1522 14520 -1470
rect 14536 -1522 14588 -1470
rect 18355 -1522 18407 -1470
rect 18423 -1522 18475 -1470
rect 18491 -1522 18543 -1470
rect 18559 -1522 18611 -1470
rect 18627 -1522 18679 -1470
rect 18695 -1522 18747 -1470
rect 18763 -1522 18815 -1470
rect 18831 -1522 18883 -1470
rect 18899 -1522 18951 -1470
rect 18967 -1522 19019 -1470
rect 19035 -1522 19087 -1470
rect 19103 -1522 19155 -1470
rect 19171 -1522 19223 -1470
rect 20196 -1522 20248 -1470
rect 20264 -1522 20316 -1470
rect 20332 -1522 20384 -1470
rect 20400 -1522 20452 -1470
rect 20468 -1522 20520 -1470
rect 20536 -1522 20588 -1470
rect 20604 -1522 20656 -1470
rect 20672 -1522 20724 -1470
rect 20740 -1522 20792 -1470
rect 20808 -1522 20860 -1470
rect 20876 -1522 20928 -1470
rect 20944 -1522 20996 -1470
rect 21012 -1522 21064 -1470
rect 6762 -7075 6814 -7023
rect 6829 -7075 6881 -7023
rect 6896 -7075 6948 -7023
rect 6963 -7075 7015 -7023
rect 7030 -7075 7082 -7023
rect 7096 -7075 7148 -7023
rect 6762 -7143 6814 -7091
rect 6829 -7143 6881 -7091
rect 6896 -7143 6948 -7091
rect 6963 -7143 7015 -7091
rect 7030 -7143 7082 -7091
rect 7096 -7143 7148 -7091
rect 3164 -7448 3216 -7396
rect 3228 -7448 3280 -7396
rect 12647 -7453 12699 -7401
rect 12739 -7453 12791 -7401
rect 12831 -7453 12883 -7401
rect 12922 -7453 12974 -7401
rect 13013 -7453 13065 -7401
rect 12647 -7557 12699 -7505
rect 12739 -7557 12791 -7505
rect 12831 -7557 12883 -7505
rect 12922 -7557 12974 -7505
rect 13013 -7557 13065 -7505
rect 8285 -7667 8337 -7615
rect 8377 -7667 8429 -7615
rect 8469 -7667 8521 -7615
rect 12647 -7661 12699 -7609
rect 12739 -7661 12791 -7609
rect 12831 -7661 12883 -7609
rect 12922 -7661 12974 -7609
rect 13013 -7661 13065 -7609
rect 5151 -8337 5203 -8285
rect 5250 -8337 5302 -8285
rect 5348 -8337 5400 -8285
rect 5151 -8411 5203 -8359
rect 5250 -8411 5302 -8359
rect 5348 -8411 5400 -8359
rect 5151 -8485 5203 -8433
rect 5250 -8485 5302 -8433
rect 5348 -8485 5400 -8433
rect 5597 -8339 5649 -8287
rect 5597 -8403 5649 -8351
rect 5597 -8467 5649 -8415
rect 5662 -8467 5906 -8287
rect 6762 -8917 6814 -8865
rect 6829 -8917 6881 -8865
rect 6896 -8917 6948 -8865
rect 6963 -8917 7015 -8865
rect 7030 -8917 7082 -8865
rect 7096 -8917 7148 -8865
rect 6762 -8985 6814 -8933
rect 6829 -8985 6881 -8933
rect 6896 -8985 6948 -8933
rect 6963 -8985 7015 -8933
rect 7030 -8985 7082 -8933
rect 7096 -8985 7148 -8933
<< metal2 >>
tri 521 16406 555 16440 ne
tri 693 16406 727 16440 nw
tri 1679 16125 1713 16159 ne
tri 1765 16125 1799 16159 nw
tri 1318 15923 1352 15957 nw
rect 803 15883 1025 15889
rect 803 15824 804 15883
rect 856 15880 888 15883
rect 940 15880 972 15883
rect 860 15824 884 15880
rect 940 15824 964 15880
rect 1024 15831 1025 15883
rect 1020 15824 1025 15831
tri 1544 15829 1578 15863 se
rect 803 15804 1025 15824
rect 803 15737 804 15804
rect 856 15793 888 15804
rect 940 15793 972 15804
rect 860 15737 884 15793
rect 940 15737 964 15793
rect 1024 15752 1025 15804
rect 1020 15737 1025 15752
rect 1402 15763 1422 15777
tri 1422 15763 1436 15777 nw
tri 1402 15743 1422 15763 nw
tri 1693 15743 1713 15763 se
rect 803 15725 1025 15737
tri 1679 15729 1693 15743 se
rect 1693 15729 1713 15743
rect 803 15650 804 15725
rect 856 15706 888 15725
rect 940 15706 972 15725
rect 860 15650 884 15706
rect 940 15650 964 15706
rect 1024 15673 1025 15725
rect 1020 15650 1025 15673
rect 803 15646 1025 15650
rect 803 15562 804 15646
rect 856 15618 888 15646
rect 940 15618 972 15646
rect 860 15562 884 15618
rect 940 15562 964 15618
rect 1024 15594 1025 15646
tri 1490 15643 1524 15677 nw
rect 1020 15588 1025 15594
rect 1020 15562 1021 15588
tri 1021 15584 1025 15588 nw
rect 803 15553 1021 15562
tri 1232 14436 1266 14470 se
tri 1320 14363 1350 14393 se
tri 1428 14311 1438 14321 se
rect 764 14281 766 14311
tri 766 14281 796 14311 nw
tri 1398 14281 1428 14311 se
rect 1428 14281 1438 14311
tri 764 14279 766 14281 nw
tri 844 14195 878 14229 nw
tri 144 12536 178 12570 nw
tri 236 11912 270 11946 nw
tri 678 8964 712 8998 se
rect 608 8894 619 8912
tri 619 8894 637 8912 nw
tri 608 8883 619 8894 nw
tri 781 8883 792 8894 se
tri 765 8867 781 8883 se
rect 781 8867 792 8883
tri 688 8786 717 8815 nw
rect 23130 7475 23270 7527
tri 23130 7445 23160 7475 ne
tri 23154 7353 23160 7359 se
rect 23160 7353 23270 7475
tri 23130 7329 23154 7353 se
rect 23154 7329 23270 7353
rect 23025 7277 23031 7329
rect 23083 7277 23097 7329
rect 23149 7277 23270 7329
tri 23130 7247 23160 7277 ne
rect 2671 7235 2692 7238
rect 2671 7186 2723 7235
rect 2671 7158 2739 7186
tri 2739 7158 2767 7186 nw
rect 2671 5387 2723 7158
tri 2723 7142 2739 7158 nw
rect 22995 7149 23051 7158
tri 23051 7128 23065 7142 sw
rect 23051 7122 23065 7128
rect 22995 7070 23013 7093
rect 22995 7069 23065 7070
rect 23051 7058 23065 7069
rect 22995 7006 23013 7013
rect 22995 7004 23065 7006
tri 23009 7000 23013 7004 ne
rect 23013 7000 23065 7004
rect 6333 6480 6339 6532
rect 6391 6529 6405 6532
rect 6457 6529 6471 6532
rect 6523 6529 6537 6532
rect 6589 6529 6603 6532
rect 6399 6480 6405 6529
rect 6655 6480 6668 6532
rect 6720 6529 6733 6532
rect 6785 6529 6798 6532
rect 6850 6529 6863 6532
rect 6915 6529 6928 6532
rect 6727 6480 6733 6529
rect 6915 6480 6917 6529
rect 6980 6480 6993 6532
rect 7045 6529 7058 6532
rect 7110 6529 7123 6532
rect 7175 6529 7188 6532
rect 7240 6529 7253 6532
rect 7055 6480 7058 6529
rect 7240 6480 7245 6529
rect 7305 6480 7318 6532
rect 7370 6529 7383 6532
rect 7435 6529 7448 6532
rect 7500 6529 7513 6532
rect 7565 6529 7578 6532
rect 7382 6480 7383 6529
rect 7565 6480 7569 6529
rect 7630 6480 7636 6532
rect 6333 6473 6343 6480
rect 6399 6473 6425 6480
rect 6481 6473 6507 6480
rect 6563 6473 6589 6480
rect 6645 6473 6671 6480
rect 6727 6473 6753 6480
rect 6809 6473 6835 6480
rect 6891 6473 6917 6480
rect 6973 6473 6999 6480
rect 7055 6473 7081 6480
rect 7137 6473 7163 6480
rect 7219 6473 7245 6480
rect 7301 6473 7326 6480
rect 7382 6473 7407 6480
rect 7463 6473 7488 6480
rect 7544 6473 7569 6480
rect 7625 6473 7636 6480
rect 6333 6421 7636 6473
rect 6333 6416 6343 6421
rect 6399 6416 6425 6421
rect 6481 6416 6507 6421
rect 6563 6416 6589 6421
rect 6645 6416 6671 6421
rect 6727 6416 6753 6421
rect 6809 6416 6835 6421
rect 6891 6416 6917 6421
rect 6973 6416 6999 6421
rect 7055 6416 7081 6421
rect 7137 6416 7163 6421
rect 7219 6416 7245 6421
rect 7301 6416 7326 6421
rect 7382 6416 7407 6421
rect 7463 6416 7488 6421
rect 7544 6416 7569 6421
rect 7625 6416 7636 6421
rect 6333 6364 6339 6416
rect 6399 6365 6405 6416
rect 6391 6364 6405 6365
rect 6457 6364 6471 6365
rect 6523 6364 6537 6365
rect 6589 6364 6603 6365
rect 6655 6364 6668 6416
rect 6727 6365 6733 6416
rect 6915 6365 6917 6416
rect 6720 6364 6733 6365
rect 6785 6364 6798 6365
rect 6850 6364 6863 6365
rect 6915 6364 6928 6365
rect 6980 6364 6993 6416
rect 7055 6365 7058 6416
rect 7240 6365 7245 6416
rect 7045 6364 7058 6365
rect 7110 6364 7123 6365
rect 7175 6364 7188 6365
rect 7240 6364 7253 6365
rect 7305 6364 7318 6416
rect 7382 6365 7383 6416
rect 7565 6365 7569 6416
rect 7370 6364 7383 6365
rect 7435 6364 7448 6365
rect 7500 6364 7513 6365
rect 7565 6364 7578 6365
rect 7630 6364 7636 6416
rect 12512 6473 12521 6529
rect 12577 6473 12606 6529
rect 12662 6473 12691 6529
rect 12747 6473 12776 6529
rect 12832 6473 12860 6529
rect 12916 6473 12944 6529
rect 13000 6473 13028 6529
rect 13084 6473 13093 6529
rect 12512 6421 13093 6473
rect 12512 6365 12521 6421
rect 12577 6365 12606 6421
rect 12662 6365 12691 6421
rect 12747 6365 12776 6421
rect 12832 6365 12860 6421
rect 12916 6365 12944 6421
rect 13000 6365 13028 6421
rect 13084 6365 13093 6421
rect 14319 6473 14328 6529
rect 14384 6473 14424 6529
rect 14480 6473 14519 6529
rect 14575 6473 14584 6529
rect 14319 6421 14584 6473
rect 14319 6365 14328 6421
rect 14384 6365 14424 6421
rect 14480 6365 14519 6421
rect 14575 6365 14584 6421
rect 18353 6480 18359 6532
rect 18411 6529 18428 6532
rect 18480 6529 18497 6532
rect 18549 6529 18565 6532
rect 18617 6529 18633 6532
rect 18685 6529 18701 6532
rect 18753 6529 18769 6532
rect 18821 6529 18837 6532
rect 18889 6529 18905 6532
rect 18957 6529 18973 6532
rect 19025 6529 19041 6532
rect 19093 6529 19109 6532
rect 19161 6529 19177 6532
rect 18419 6480 18428 6529
rect 18685 6480 18687 6529
rect 18753 6480 18768 6529
rect 18824 6480 18837 6529
rect 19161 6480 19169 6529
rect 19229 6480 19235 6532
rect 18353 6473 18363 6480
rect 18419 6473 18444 6480
rect 18500 6473 18525 6480
rect 18581 6473 18606 6480
rect 18662 6473 18687 6480
rect 18743 6473 18768 6480
rect 18824 6473 18849 6480
rect 18905 6473 18929 6480
rect 18985 6473 19009 6480
rect 19065 6473 19089 6480
rect 19145 6473 19169 6480
rect 19225 6473 19235 6480
rect 18353 6421 19235 6473
rect 18353 6416 18363 6421
rect 18419 6416 18444 6421
rect 18500 6416 18525 6421
rect 18581 6416 18606 6421
rect 18662 6416 18687 6421
rect 18743 6416 18768 6421
rect 18824 6416 18849 6421
rect 18905 6416 18929 6421
rect 18985 6416 19009 6421
rect 19065 6416 19089 6421
rect 19145 6416 19169 6421
rect 19225 6416 19235 6421
rect 18353 6364 18359 6416
rect 18419 6365 18428 6416
rect 18685 6365 18687 6416
rect 18753 6365 18768 6416
rect 18824 6365 18837 6416
rect 19161 6365 19169 6416
rect 18411 6364 18428 6365
rect 18480 6364 18497 6365
rect 18549 6364 18565 6365
rect 18617 6364 18633 6365
rect 18685 6364 18701 6365
rect 18753 6364 18769 6365
rect 18821 6364 18837 6365
rect 18889 6364 18905 6365
rect 18957 6364 18973 6365
rect 19025 6364 19041 6365
rect 19093 6364 19109 6365
rect 19161 6364 19177 6365
rect 19229 6364 19235 6416
rect 20192 6480 20198 6532
rect 20250 6529 20267 6532
rect 20319 6529 20336 6532
rect 20388 6529 20404 6532
rect 20456 6529 20472 6532
rect 20524 6529 20540 6532
rect 20592 6529 20608 6532
rect 20660 6529 20676 6532
rect 20728 6529 20744 6532
rect 20796 6529 20812 6532
rect 20864 6529 20880 6532
rect 20932 6529 20948 6532
rect 21000 6529 21016 6532
rect 20258 6480 20267 6529
rect 20524 6480 20526 6529
rect 20592 6480 20607 6529
rect 20663 6480 20676 6529
rect 21000 6480 21008 6529
rect 21068 6480 21074 6532
rect 20192 6473 20202 6480
rect 20258 6473 20283 6480
rect 20339 6473 20364 6480
rect 20420 6473 20445 6480
rect 20501 6473 20526 6480
rect 20582 6473 20607 6480
rect 20663 6473 20688 6480
rect 20744 6473 20768 6480
rect 20824 6473 20848 6480
rect 20904 6473 20928 6480
rect 20984 6473 21008 6480
rect 21064 6473 21074 6480
rect 20192 6421 21074 6473
rect 20192 6416 20202 6421
rect 20258 6416 20283 6421
rect 20339 6416 20364 6421
rect 20420 6416 20445 6421
rect 20501 6416 20526 6421
rect 20582 6416 20607 6421
rect 20663 6416 20688 6421
rect 20744 6416 20768 6421
rect 20824 6416 20848 6421
rect 20904 6416 20928 6421
rect 20984 6416 21008 6421
rect 21064 6416 21074 6421
rect 20192 6364 20198 6416
rect 20258 6365 20267 6416
rect 20524 6365 20526 6416
rect 20592 6365 20607 6416
rect 20663 6365 20676 6416
rect 21000 6365 21008 6416
rect 20250 6364 20267 6365
rect 20319 6364 20336 6365
rect 20388 6364 20404 6365
rect 20456 6364 20472 6365
rect 20524 6364 20540 6365
rect 20592 6364 20608 6365
rect 20660 6364 20676 6365
rect 20728 6364 20744 6365
rect 20796 6364 20812 6365
rect 20864 6364 20880 6365
rect 20932 6364 20948 6365
rect 21000 6364 21016 6365
rect 21068 6364 21074 6416
rect 22975 6480 22981 6532
rect 23033 6529 23072 6532
rect 22975 6473 22985 6480
rect 23041 6473 23065 6529
rect 23124 6480 23130 6532
rect 23121 6473 23130 6480
rect 22975 6421 23130 6473
rect 22975 6416 22985 6421
rect 22975 6364 22981 6416
rect 23041 6365 23065 6421
rect 23121 6416 23130 6421
rect 23033 6364 23072 6365
rect 23124 6364 23130 6416
tri 23154 5779 23160 5785 se
rect 23160 5779 23270 7277
rect 25109 7353 25916 7359
rect 25225 7311 25916 7353
tri 25916 7311 25964 7359 sw
rect 25225 7237 25964 7311
rect 25109 7231 25964 7237
tri 25795 7183 25843 7231 ne
rect 25105 7122 25673 7128
rect 25221 7080 25673 7122
tri 25673 7080 25721 7128 sw
rect 25221 7006 25721 7080
rect 25105 7000 25721 7006
tri 25537 6967 25570 7000 ne
rect 23154 5773 23270 5779
rect 23154 5587 23270 5593
rect 8088 5550 8216 5552
rect 8088 5498 8094 5550
rect 8146 5498 8158 5550
rect 8210 5498 8216 5550
tri 2723 5387 2725 5389 sw
rect 6121 5387 6127 5439
rect 6179 5387 6191 5439
rect 6243 5387 6249 5439
rect 2671 5364 2725 5387
tri 2725 5364 2748 5387 sw
rect 2671 5320 2961 5364
rect 2671 5312 2740 5320
tri 2740 5312 2748 5320 nw
tri 2902 5312 2910 5320 ne
rect 2910 5312 2961 5320
rect 2963 5312 3041 5364
rect 3093 5312 3105 5364
rect 3157 5312 3163 5364
rect 2435 5190 2441 5242
rect 2493 5190 2505 5242
rect 2557 5190 2563 5242
rect 2508 5103 2514 5155
rect 2566 5103 2578 5155
rect 2630 5103 2636 5155
rect 2671 5070 2723 5312
tri 2723 5295 2740 5312 nw
tri 6111 5217 6121 5227 se
rect 6121 5217 6249 5387
tri 6089 5195 6111 5217 se
rect 6111 5195 6249 5217
tri 5479 5177 5497 5195 se
rect 5497 5177 6249 5195
tri 5467 5165 5479 5177 se
rect 5479 5165 6249 5177
tri 6249 5165 6261 5177 sw
tri 5466 5164 5467 5165 se
rect 5467 5164 6261 5165
rect 5466 5142 6261 5164
tri 6261 5142 6284 5165 sw
rect 5466 5120 6380 5142
tri 6380 5120 6402 5142 sw
rect 5466 5116 6402 5120
rect 5466 5105 5633 5116
tri 5633 5105 5644 5116 nw
tri 6176 5105 6187 5116 ne
rect 6187 5105 6402 5116
tri 2723 5070 2758 5105 sw
tri 5449 4966 5466 4983 se
rect 5466 4966 5618 5105
tri 5618 5090 5633 5105 nw
tri 6187 5090 6202 5105 ne
rect 6202 5090 6402 5105
tri 6202 5070 6222 5090 ne
rect 6222 5070 6402 5090
tri 6222 5018 6274 5070 ne
rect 6274 5018 6402 5070
rect 8088 5018 8202 5498
tri 8202 5484 8216 5498 nw
rect 11308 5550 11436 5552
rect 11308 5498 11314 5550
rect 11366 5498 11378 5550
rect 11430 5498 11436 5550
tri 8202 5018 8248 5064 sw
rect 11308 5018 11422 5498
tri 11422 5484 11436 5498 nw
rect 14528 5550 14656 5552
rect 14528 5498 14534 5550
rect 14586 5498 14598 5550
rect 14650 5498 14656 5550
tri 13290 5064 13293 5067 se
rect 13293 5064 13823 5067
tri 13823 5064 13826 5067 sw
tri 11422 5018 11468 5064 sw
tri 13244 5018 13290 5064 se
rect 13290 5018 13826 5064
tri 13826 5018 13872 5064 sw
rect 14528 5018 14642 5498
tri 14642 5484 14656 5498 nw
rect 17748 5550 17876 5552
rect 17748 5498 17754 5550
rect 17806 5498 17818 5550
rect 17870 5498 17876 5550
rect 16264 5165 16270 5217
rect 16322 5165 16337 5217
rect 16389 5165 16404 5217
rect 16456 5165 16470 5217
rect 16522 5165 16528 5217
tri 14642 5018 14688 5064 sw
rect 6274 4966 6280 5018
rect 6332 4966 6344 5018
rect 6396 4966 6402 5018
rect 7632 4966 7638 5018
rect 7690 4966 7702 5018
rect 7754 5005 7780 5018
tri 7780 5005 7793 5018 sw
rect 7754 4966 7793 5005
tri 5436 4953 5449 4966 se
rect 5449 4953 5618 4966
tri 7720 4965 7721 4966 ne
rect 7721 4965 7793 4966
tri 5618 4953 5630 4965 sw
tri 7721 4953 7733 4965 ne
tri 5423 4940 5436 4953 se
rect 5436 4940 5630 4953
tri 5630 4940 5643 4953 sw
rect 5423 4888 5429 4940
rect 5481 4888 5507 4940
rect 5559 4888 5585 4940
rect 5637 4888 5643 4940
rect 2680 4734 2686 4786
rect 2738 4734 2750 4786
rect 2802 4734 2808 4786
rect 7733 4400 7793 4965
tri 13213 4987 13244 5018 se
rect 13244 4987 13872 5018
rect 13213 4983 13872 4987
tri 13872 4983 13907 5018 sw
rect 13213 4940 13349 4983
tri 13349 4940 13392 4983 nw
tri 13722 4940 13765 4983 ne
rect 13765 4981 13907 4983
tri 13907 4981 13909 4983 sw
rect 13765 4940 13909 4981
rect 7833 4888 7839 4940
rect 7891 4888 7908 4940
rect 7960 4888 7976 4940
rect 8028 4888 8034 4940
rect 7833 4506 8034 4888
rect 8692 4506 8820 4792
rect 7833 4454 7839 4506
rect 7891 4454 7908 4506
rect 7960 4454 7976 4506
rect 8028 4454 8034 4506
rect 8086 4454 8092 4506
rect 8144 4454 8156 4506
rect 8208 4454 8214 4506
rect 8692 4454 8698 4506
rect 8750 4454 8762 4506
rect 8814 4454 8820 4506
rect 11912 4506 12040 4792
rect 11912 4454 11918 4506
rect 11970 4454 11982 4506
rect 12034 4454 12040 4506
rect 13213 4506 13341 4940
tri 13341 4932 13349 4940 nw
rect 13213 4454 13219 4506
rect 13271 4454 13283 4506
rect 13335 4454 13341 4506
rect 13444 4888 13450 4940
rect 13502 4888 13519 4940
rect 13571 4888 13587 4940
rect 13639 4888 13645 4940
tri 13765 4932 13773 4940 ne
rect 13773 4932 13909 4940
tri 13773 4924 13781 4932 ne
rect 8086 4444 8159 4454
tri 8159 4444 8169 4454 nw
rect 13444 4444 13645 4888
rect 13781 4506 13909 4932
rect 16264 4940 16528 5165
rect 17748 5018 17862 5498
tri 17862 5484 17876 5498 nw
rect 20968 5550 21096 5552
rect 20968 5498 20974 5550
rect 21026 5498 21038 5550
rect 21090 5498 21096 5550
tri 19370 5064 19373 5067 se
rect 19373 5064 19903 5067
tri 19903 5064 19906 5067 sw
tri 17862 5018 17908 5064 sw
tri 19324 5018 19370 5064 se
rect 19370 5018 19906 5064
tri 19906 5018 19952 5064 sw
rect 20968 5018 21082 5498
tri 21082 5484 21096 5498 nw
rect 24188 5550 24316 5552
rect 24188 5498 24194 5550
rect 24246 5498 24258 5550
rect 24310 5498 24316 5550
rect 23347 5166 23353 5282
rect 23469 5166 23475 5282
tri 23288 5067 23347 5126 se
rect 23347 5069 23475 5166
rect 23347 5067 23473 5069
tri 23473 5067 23475 5069 nw
tri 22707 5064 22710 5067 se
rect 22710 5064 23424 5067
tri 21082 5018 21128 5064 sw
tri 22661 5018 22707 5064 se
rect 22707 5018 23424 5064
tri 23424 5018 23473 5067 nw
rect 24188 5018 24302 5498
tri 24302 5484 24316 5498 nw
rect 25570 5439 25721 7000
rect 25570 5323 25583 5439
rect 25699 5323 25721 5439
rect 24792 5266 24920 5282
rect 24792 5214 24798 5266
rect 24850 5214 24862 5266
rect 24914 5214 24920 5266
tri 24302 5018 24348 5064 sw
tri 24749 5018 24792 5061 se
rect 24792 5018 24920 5214
tri 24920 5018 24963 5061 sw
rect 16264 4888 16270 4940
rect 16322 4888 16337 4940
rect 16389 4888 16404 4940
rect 16456 4888 16470 4940
rect 16522 4888 16528 4940
tri 19293 4987 19324 5018 se
rect 19324 4987 19952 5018
rect 19293 4983 19952 4987
tri 19952 4983 19987 5018 sw
tri 22630 4987 22661 5018 se
rect 22661 4987 23393 5018
tri 23393 4987 23424 5018 nw
rect 22630 4983 23389 4987
tri 23389 4983 23393 4987 nw
rect 19293 4940 19429 4983
tri 19429 4940 19472 4983 nw
tri 19802 4940 19845 4983 ne
rect 19845 4981 19987 4983
tri 19987 4981 19989 4983 sw
rect 19845 4940 19989 4981
rect 13781 4454 13787 4506
rect 13839 4454 13851 4506
rect 13903 4454 13909 4506
rect 15132 4506 15260 4792
rect 15132 4454 15138 4506
rect 15190 4454 15202 4506
rect 15254 4454 15260 4506
rect 18352 4506 18480 4792
rect 18352 4454 18358 4506
rect 18410 4454 18422 4506
rect 18474 4454 18480 4506
rect 19293 4506 19421 4940
tri 19421 4932 19429 4940 nw
rect 19513 4888 19519 4940
rect 19571 4888 19588 4940
rect 19640 4888 19656 4940
rect 19708 4888 19714 4940
tri 19845 4932 19853 4940 ne
rect 19853 4932 19989 4940
tri 19853 4924 19861 4932 ne
rect 19513 4566 19714 4888
rect 19513 4514 19519 4566
rect 19571 4514 19588 4566
rect 19640 4514 19656 4566
rect 19708 4514 19714 4566
rect 19293 4454 19299 4506
rect 19351 4454 19363 4506
rect 19415 4454 19421 4506
rect 19861 4506 19989 4932
rect 22630 4940 22766 4983
tri 22766 4940 22809 4983 nw
rect 19861 4454 19867 4506
rect 19919 4454 19931 4506
rect 19983 4454 19989 4506
rect 21572 4506 21700 4792
rect 21572 4454 21578 4506
rect 21630 4454 21642 4506
rect 21694 4454 21700 4506
rect 22630 4506 22758 4940
tri 22758 4932 22766 4940 nw
rect 22907 4888 22913 4940
rect 22965 4888 22982 4940
rect 23034 4888 23050 4940
rect 23102 4888 23108 4940
rect 22907 4626 23108 4888
rect 22907 4574 22913 4626
rect 22965 4574 22982 4626
rect 23034 4574 23050 4626
rect 23102 4574 23108 4626
rect 25570 4660 25721 5323
tri 25811 5288 25843 5320 se
rect 25843 5288 25964 7231
rect 26101 5338 26107 5360
tri 26101 5332 26107 5338 ne
tri 26107 5332 26135 5360 nw
rect 25789 5282 25964 5288
rect 25789 5166 25842 5282
rect 25958 5166 25964 5282
rect 25789 5160 25964 5166
tri 25721 4660 25795 4734 sw
rect 22630 4454 22636 4506
rect 22688 4454 22700 4506
rect 22752 4454 22758 4506
rect 23657 4500 23663 4616
rect 23779 4500 23785 4616
rect 25570 4544 25742 4660
rect 25858 4544 25864 4660
tri 25983 4461 25986 4464 se
tri 26034 4457 26038 4461 nw
rect 8086 4440 8155 4444
tri 8155 4440 8159 4444 nw
tri 8081 4435 8086 4440 se
rect 8086 4435 8115 4440
tri 7793 4400 7828 4435 sw
tri 8046 4400 8081 4435 se
rect 8081 4400 8115 4435
tri 8115 4400 8155 4440 nw
rect 7733 4392 8107 4400
tri 8107 4392 8115 4400 nw
rect 13444 4392 13450 4444
rect 13502 4392 13519 4444
rect 13571 4392 13587 4444
rect 13639 4392 13645 4444
rect 7733 4391 8106 4392
tri 8106 4391 8107 4392 nw
tri 7733 4353 7771 4391 ne
rect 7771 4353 8068 4391
tri 8068 4353 8106 4391 nw
rect 23472 4082 23623 4120
rect 8386 3591 8803 3697
rect 2844 2470 2896 2476
rect 2844 2406 2896 2418
rect 2326 1758 2378 1764
tri 2296 1706 2315 1725 ne
rect 2315 1706 2326 1725
tri 2315 1695 2326 1706 ne
rect 2326 1694 2378 1706
tri 2215 1637 2219 1641 ne
rect 2219 1637 2242 1641
tri 512 1609 540 1637 sw
tri 2219 1614 2242 1637 ne
rect 2326 1636 2378 1642
rect 2844 1758 2896 2354
rect 2995 2470 3047 3365
tri 20185 3083 20189 3087 se
tri 20185 2889 20189 2893 ne
rect 2995 2406 3047 2418
rect 2995 2348 3047 2354
tri 20976 2259 20980 2263 se
rect 20980 2259 20983 2263
tri 20976 2065 20980 2069 ne
rect 20980 2065 20983 2069
rect 2844 1694 2896 1706
rect 2844 1636 2896 1642
tri 2131 1553 2135 1557 ne
rect 2135 1553 2158 1557
tri 420 1525 448 1553 sw
tri 2135 1530 2158 1553 ne
tri 2044 1469 2048 1473 ne
rect 2048 1469 2074 1473
tri 328 1441 356 1469 sw
tri 2048 1443 2074 1469 ne
tri 1961 1385 1965 1389 ne
rect 1965 1385 1990 1389
tri 236 1357 264 1385 sw
tri 1965 1360 1990 1385 ne
rect 24034 1346 24912 2591
tri 1875 1301 1879 1305 ne
rect 1879 1301 1906 1305
tri 144 1286 159 1301 sw
tri 1879 1286 1894 1301 ne
rect 1894 1286 1906 1301
rect 144 1280 159 1286
tri 159 1280 165 1286 sw
tri 1894 1280 1900 1286 ne
rect 1900 1280 1906 1286
rect 144 1273 165 1280
tri 165 1273 172 1280 sw
tri 1900 1274 1906 1280 ne
rect 23704 1280 23789 1292
rect 23704 1228 23720 1280
rect 23772 1228 23789 1280
tri 1796 1217 1800 1221 ne
rect 1800 1217 1822 1221
tri 52 1216 53 1217 sw
tri 1800 1216 1801 1217 ne
rect 1801 1216 1822 1217
rect 52 1189 53 1216
tri 53 1189 80 1216 sw
tri 1801 1195 1822 1216 ne
rect 23704 1216 23789 1228
rect 23704 1164 23720 1216
rect 23772 1164 23789 1216
rect 23704 1152 23789 1164
tri 1708 1107 1738 1137 ne
rect 23704 1100 23720 1152
rect 23772 1100 23789 1152
tri 26468 1111 26502 1145 ne
rect 2004 765 2031 792
tri 2241 -376 2326 -291 se
rect 2326 -324 2378 947
tri 3684 812 3718 846 ne
tri 2896 748 2930 782 sw
rect 2844 696 2850 748
rect 2902 696 2914 748
rect 2966 696 2972 748
tri 2896 662 2930 696 nw
tri 6836 577 6838 579 se
tri 3141 494 3171 524 sw
tri 9316 500 9318 502 se
tri 9721 500 9723 502 sw
tri 10247 500 10249 502 se
tri 10249 500 10251 502 sw
tri 10650 500 10652 502 se
tri 10652 500 10654 502 sw
tri 15804 500 15806 502 se
tri 16209 500 16211 502 sw
tri 16731 500 16733 502 se
tri 17136 500 17138 502 sw
tri 22369 500 22371 502 se
tri 22693 500 22695 502 sw
tri 10246 499 10247 500 se
rect 10247 499 10251 500
tri 10251 499 10252 500 sw
tri 10649 499 10650 500 se
rect 10650 499 10654 500
tri 10654 499 10655 500 sw
rect 3141 490 3171 494
tri 3171 490 3175 494 sw
tri 3614 490 3618 494 sw
rect 3614 449 3618 490
tri 3618 449 3659 490 sw
tri 10246 448 10247 449 ne
rect 10247 448 10249 449
tri 9316 446 9318 448 ne
tri 9721 446 9723 448 nw
tri 10247 446 10249 448 ne
tri 10249 446 10252 449 nw
tri 10649 446 10652 449 ne
tri 10652 446 10655 449 nw
tri 15803 446 15806 449 ne
tri 16209 446 16212 449 nw
tri 16730 446 16733 449 ne
tri 17136 446 17139 449 nw
tri 22368 446 22371 449 ne
tri 22693 446 22696 449 nw
tri 3141 404 3175 438 nw
tri 6889 374 6910 395 sw
tri 6823 361 6836 374 se
rect 6889 361 6910 374
tri 6910 361 6923 374 sw
tri 9316 188 9318 190 se
tri 9721 188 9723 190 sw
tri 10247 188 10249 190 se
tri 10249 188 10251 190 sw
tri 10650 188 10652 190 se
tri 10652 188 10654 190 sw
tri 15800 188 15802 190 se
tri 16205 188 16207 190 sw
tri 16731 188 16733 190 se
tri 17136 188 17138 190 sw
tri 22369 188 22371 190 se
tri 22689 188 22691 190 sw
tri 10246 187 10247 188 se
rect 10247 187 10251 188
tri 10251 187 10252 188 sw
tri 10649 187 10650 188 se
rect 10650 187 10654 188
tri 10654 187 10655 188 sw
tri 10246 136 10247 137 ne
rect 10247 136 10249 137
tri 9316 134 9318 136 ne
tri 9721 134 9723 136 nw
tri 10247 134 10249 136 ne
tri 10249 134 10252 137 nw
tri 10649 134 10652 137 ne
tri 10652 134 10655 137 nw
tri 15799 134 15802 137 ne
tri 16205 134 16208 137 nw
tri 16730 134 16733 137 ne
tri 17136 134 17139 137 nw
tri 22368 134 22371 137 ne
tri 22689 134 22692 137 nw
rect 2844 -72 2850 -20
rect 2902 -72 2914 -20
rect 2966 -72 2972 -20
tri 9316 -124 9318 -122 se
tri 9721 -124 9723 -122 sw
tri 10247 -124 10249 -122 se
tri 10249 -124 10251 -122 sw
tri 10650 -124 10652 -122 se
tri 10652 -124 10654 -122 sw
tri 15800 -124 15802 -122 se
tri 16205 -124 16207 -122 sw
tri 16731 -124 16733 -122 se
tri 17136 -124 17138 -122 sw
tri 22369 -124 22371 -122 se
tri 22689 -124 22691 -122 sw
tri 10246 -125 10247 -124 se
rect 10247 -125 10251 -124
tri 10251 -125 10252 -124 sw
tri 10649 -125 10650 -124 se
rect 10650 -125 10654 -124
tri 10654 -125 10655 -124 sw
tri 10246 -176 10247 -175 ne
rect 10247 -176 10249 -175
tri 9316 -178 9318 -176 ne
tri 9721 -178 9723 -176 nw
tri 10247 -178 10249 -176 ne
tri 10249 -178 10252 -175 nw
tri 10649 -178 10652 -175 ne
tri 10652 -178 10655 -175 nw
tri 15799 -178 15802 -175 ne
tri 16205 -178 16208 -175 nw
tri 16730 -178 16733 -175 ne
tri 17136 -178 17139 -175 nw
tri 22368 -178 22371 -175 ne
tri 22689 -178 22692 -175 nw
tri 2326 -376 2378 -324 nw
tri 2229 -388 2241 -376 se
rect 2241 -388 2314 -376
tri 2314 -388 2326 -376 nw
tri 2204 -481 2229 -456 se
rect 2229 -481 2285 -388
tri 2285 -417 2314 -388 nw
rect 23704 -417 23789 1100
tri 23789 -417 23796 -410 sw
rect 23704 -418 23796 -417
tri 23796 -418 23797 -417 sw
rect 23704 -423 23797 -418
tri 23797 -423 23802 -418 sw
tri 25703 -423 25708 -418 nw
rect 2157 -533 2163 -481
rect 2215 -533 2227 -481
rect 2279 -533 2285 -481
tri 23668 -481 23704 -445 se
rect 23704 -481 23802 -423
tri 23802 -481 23860 -423 sw
rect 23668 -533 23674 -481
rect 23726 -533 23738 -481
rect 23790 -533 23802 -481
rect 23854 -533 23860 -481
rect 13711 -1459 13720 -1403
rect 13776 -1459 13801 -1403
rect 13857 -1459 13882 -1403
rect 13938 -1459 13963 -1403
rect 14019 -1459 14044 -1403
rect 14100 -1459 14125 -1403
rect 14181 -1459 14206 -1403
rect 14262 -1459 14286 -1403
rect 14342 -1459 14366 -1403
rect 14422 -1459 14446 -1403
rect 14502 -1459 14526 -1403
rect 14582 -1459 14594 -1403
rect 13711 -1470 14594 -1459
rect 13711 -1522 13720 -1470
rect 13772 -1522 13788 -1470
rect 13840 -1522 13856 -1470
rect 13908 -1522 13924 -1470
rect 13976 -1522 13992 -1470
rect 14044 -1522 14060 -1470
rect 14112 -1522 14128 -1470
rect 14180 -1522 14196 -1470
rect 14248 -1522 14264 -1470
rect 14316 -1522 14332 -1470
rect 14384 -1522 14400 -1470
rect 14452 -1522 14468 -1470
rect 14520 -1522 14536 -1470
rect 14588 -1522 14594 -1470
rect 18349 -1409 18358 -1353
rect 18414 -1409 18439 -1353
rect 18495 -1409 18520 -1353
rect 18576 -1409 18601 -1353
rect 18657 -1409 18682 -1353
rect 18738 -1409 18763 -1353
rect 18819 -1409 18844 -1353
rect 18900 -1409 18924 -1353
rect 18980 -1409 19004 -1353
rect 19060 -1409 19084 -1353
rect 19140 -1409 19164 -1353
rect 19220 -1409 19229 -1353
rect 18349 -1461 19229 -1409
rect 18349 -1470 18358 -1461
rect 18414 -1470 18439 -1461
rect 18495 -1470 18520 -1461
rect 18576 -1470 18601 -1461
rect 18657 -1470 18682 -1461
rect 18738 -1470 18763 -1461
rect 18819 -1470 18844 -1461
rect 18900 -1470 18924 -1461
rect 18980 -1470 19004 -1461
rect 19060 -1470 19084 -1461
rect 19140 -1470 19164 -1461
rect 19220 -1470 19229 -1461
rect 18349 -1522 18355 -1470
rect 18414 -1517 18423 -1470
rect 18679 -1517 18682 -1470
rect 18407 -1522 18423 -1517
rect 18475 -1522 18491 -1517
rect 18543 -1522 18559 -1517
rect 18611 -1522 18627 -1517
rect 18679 -1522 18695 -1517
rect 18747 -1522 18763 -1470
rect 18819 -1517 18831 -1470
rect 19155 -1517 19164 -1470
rect 18815 -1522 18831 -1517
rect 18883 -1522 18899 -1517
rect 18951 -1522 18967 -1517
rect 19019 -1522 19035 -1517
rect 19087 -1522 19103 -1517
rect 19155 -1522 19171 -1517
rect 19223 -1522 19229 -1470
rect 20190 -1409 20199 -1353
rect 20255 -1409 20280 -1353
rect 20336 -1409 20361 -1353
rect 20417 -1409 20442 -1353
rect 20498 -1409 20523 -1353
rect 20579 -1409 20604 -1353
rect 20660 -1409 20685 -1353
rect 20741 -1409 20765 -1353
rect 20821 -1409 20845 -1353
rect 20901 -1409 20925 -1353
rect 20981 -1409 21005 -1353
rect 21061 -1409 21070 -1353
rect 20190 -1461 21070 -1409
rect 20190 -1470 20199 -1461
rect 20255 -1470 20280 -1461
rect 20336 -1470 20361 -1461
rect 20417 -1470 20442 -1461
rect 20498 -1470 20523 -1461
rect 20579 -1470 20604 -1461
rect 20660 -1470 20685 -1461
rect 20741 -1470 20765 -1461
rect 20821 -1470 20845 -1461
rect 20901 -1470 20925 -1461
rect 20981 -1470 21005 -1461
rect 21061 -1470 21070 -1461
rect 20190 -1522 20196 -1470
rect 20255 -1517 20264 -1470
rect 20520 -1517 20523 -1470
rect 20248 -1522 20264 -1517
rect 20316 -1522 20332 -1517
rect 20384 -1522 20400 -1517
rect 20452 -1522 20468 -1517
rect 20520 -1522 20536 -1517
rect 20588 -1522 20604 -1470
rect 20660 -1517 20672 -1470
rect 20996 -1517 21005 -1470
rect 20656 -1522 20672 -1517
rect 20724 -1522 20740 -1517
rect 20792 -1522 20808 -1517
rect 20860 -1522 20876 -1517
rect 20928 -1522 20944 -1517
rect 20996 -1522 21012 -1517
rect 21064 -1522 21070 -1470
rect 26647 -5487 26930 -5417
tri 26574 -6180 26608 -6146 se
rect 6756 -7075 6762 -7023
rect 6814 -7056 6829 -7023
rect 6881 -7056 6896 -7023
rect 6948 -7056 6963 -7023
rect 7015 -7056 7030 -7023
rect 7082 -7056 7096 -7023
rect 6822 -7075 6829 -7056
rect 7082 -7075 7088 -7056
rect 7148 -7075 7154 -7023
rect 6756 -7091 6766 -7075
rect 6822 -7091 6847 -7075
rect 6903 -7091 6928 -7075
rect 6984 -7091 7008 -7075
rect 7064 -7091 7088 -7075
rect 7144 -7091 7154 -7075
rect 6756 -7143 6762 -7091
rect 6822 -7112 6829 -7091
rect 7082 -7112 7088 -7091
rect 6814 -7143 6829 -7112
rect 6881 -7143 6896 -7112
rect 6948 -7143 6963 -7112
rect 7015 -7143 7030 -7112
rect 7082 -7143 7096 -7112
rect 7148 -7143 7154 -7091
tri 6488 -7361 6509 -7340 ne
rect 6509 -7361 6522 -7340
tri 3162 -7366 3167 -7361 se
rect 3167 -7366 3223 -7361
tri 3223 -7366 3228 -7361 sw
tri 6509 -7366 6514 -7361 ne
rect 6514 -7366 6522 -7361
rect 3158 -7370 3260 -7366
rect 3158 -7396 3167 -7370
rect 3223 -7396 3260 -7370
tri 6514 -7374 6522 -7366 ne
rect 3158 -7448 3164 -7396
rect 3223 -7426 3228 -7396
rect 3216 -7448 3228 -7426
rect 3280 -7448 3286 -7396
rect 12636 -7399 13078 -7398
tri 3158 -7453 3163 -7448 ne
rect 3163 -7450 3252 -7448
rect 3163 -7453 3167 -7450
tri 3163 -7457 3167 -7453 ne
rect 3223 -7453 3252 -7450
tri 3252 -7453 3257 -7448 nw
rect 3223 -7457 3248 -7453
tri 3248 -7457 3252 -7453 nw
rect 12636 -7455 12645 -7399
rect 12701 -7401 12768 -7399
rect 12824 -7401 12891 -7399
rect 12947 -7401 13013 -7399
rect 12701 -7453 12739 -7401
rect 12824 -7453 12831 -7401
rect 12883 -7453 12891 -7401
rect 12974 -7453 13013 -7401
rect 12701 -7455 12768 -7453
rect 12824 -7455 12891 -7453
rect 12947 -7455 13013 -7453
rect 13069 -7455 13078 -7399
tri 3223 -7482 3248 -7457 nw
rect 3167 -7515 3223 -7506
rect 12636 -7503 13078 -7455
rect 12636 -7559 12645 -7503
rect 12701 -7505 12768 -7503
rect 12824 -7505 12891 -7503
rect 12947 -7505 13013 -7503
rect 12701 -7557 12739 -7505
rect 12824 -7557 12831 -7505
rect 12883 -7557 12891 -7505
rect 12974 -7557 13013 -7505
rect 12701 -7559 12768 -7557
rect 12824 -7559 12891 -7557
rect 12947 -7559 13013 -7557
rect 13069 -7559 13078 -7503
rect 12636 -7607 13078 -7559
rect 8265 -7669 8274 -7613
rect 8330 -7615 8371 -7613
rect 8427 -7615 8467 -7613
rect 8337 -7667 8371 -7615
rect 8429 -7667 8467 -7615
rect 8330 -7669 8371 -7667
rect 8427 -7669 8467 -7667
rect 8523 -7669 8532 -7613
rect 12636 -7663 12645 -7607
rect 12701 -7609 12768 -7607
rect 12824 -7609 12891 -7607
rect 12947 -7609 13013 -7607
rect 12701 -7661 12739 -7609
rect 12824 -7661 12831 -7609
rect 12883 -7661 12891 -7609
rect 12974 -7661 13013 -7609
rect 12701 -7663 12768 -7661
rect 12824 -7663 12891 -7661
rect 12947 -7663 13013 -7661
rect 13069 -7663 13078 -7607
rect 12636 -7664 13078 -7663
tri 1669 -7733 1697 -7705 ne
rect 1697 -7733 1703 -7705
tri 1743 -7733 1771 -7705 nw
tri 1697 -7739 1703 -7733 ne
tri 11162 -7782 11174 -7770 se
tri 8340 -7820 8352 -7808 ne
rect 8352 -7820 8353 -7808
tri 8976 -7894 9010 -7860 ne
rect 9010 -7894 9014 -7860
tri 9010 -7898 9014 -7894 ne
tri 11218 -7898 11222 -7894 ne
rect 11222 -7898 11238 -7894
tri 11222 -7907 11231 -7898 ne
rect 11231 -7907 11238 -7898
rect 8469 -7928 8470 -7921
tri 8470 -7928 8477 -7921 sw
rect 8465 -7973 8470 -7962
tri 8470 -7973 8481 -7962 nw
tri 5577 -8008 5587 -7998 sw
tri 768 -8011 771 -8008 sw
rect 5576 -8048 5579 -8008
rect 5576 -8050 5577 -8048
tri 5577 -8050 5579 -8048 nw
tri 11967 -8067 11983 -8051 ne
rect 11983 -8067 11990 -8051
tri 769 -8137 771 -8135 nw
tri 8571 -8196 8584 -8183 se
rect 8584 -8196 8585 -8183
tri 8550 -8270 8579 -8241 ne
rect 8579 -8270 8584 -8241
rect 5132 -8326 5141 -8270
rect 5197 -8285 5252 -8270
rect 5308 -8285 5363 -8270
rect 5132 -8337 5151 -8326
rect 5203 -8337 5250 -8285
rect 5308 -8326 5348 -8285
rect 5419 -8326 5428 -8270
tri 8579 -8275 8584 -8270 ne
rect 5302 -8337 5348 -8326
rect 5400 -8337 5428 -8326
rect 5132 -8354 5428 -8337
rect 5132 -8410 5141 -8354
rect 5197 -8359 5252 -8354
rect 5308 -8359 5363 -8354
rect 5132 -8411 5151 -8410
rect 5203 -8411 5250 -8359
rect 5308 -8410 5348 -8359
rect 5419 -8410 5428 -8354
rect 5302 -8411 5348 -8410
rect 5400 -8411 5428 -8410
rect 5132 -8433 5428 -8411
rect 5132 -8438 5151 -8433
rect 5132 -8494 5141 -8438
rect 5203 -8485 5250 -8433
rect 5302 -8438 5348 -8433
rect 5400 -8438 5428 -8433
rect 5308 -8485 5348 -8438
rect 5197 -8494 5252 -8485
rect 5308 -8494 5363 -8485
rect 5419 -8494 5428 -8438
rect 5584 -8343 5593 -8287
rect 5649 -8343 5662 -8287
rect 5912 -8343 5921 -8287
tri 12339 -8290 12340 -8289 ne
rect 12340 -8290 12362 -8289
tri 8334 -8305 8349 -8290 se
rect 8349 -8299 8455 -8290
rect 8349 -8305 8374 -8299
tri 8331 -8308 8334 -8305 se
rect 8334 -8308 8374 -8305
rect 5584 -8351 5662 -8343
rect 5584 -8403 5597 -8351
rect 5649 -8403 5662 -8351
rect 5584 -8411 5662 -8403
rect 5906 -8411 5921 -8343
rect 8317 -8355 8374 -8308
rect 8430 -8355 8455 -8299
tri 12340 -8305 12355 -8290 ne
rect 12355 -8305 12362 -8290
rect 8317 -8360 8455 -8355
tri 8317 -8387 8344 -8360 ne
rect 8344 -8379 8455 -8360
rect 5584 -8467 5593 -8411
rect 5649 -8467 5662 -8411
rect 5912 -8467 5921 -8411
rect 8344 -8435 8374 -8379
rect 8430 -8435 8455 -8379
rect 8344 -8444 8455 -8435
tri 6402 -8676 6404 -8674 nw
rect 3425 -8842 3430 -8833
tri 3430 -8842 3439 -8833 sw
rect 3425 -8854 3439 -8842
tri 3439 -8854 3451 -8842 sw
tri 13151 -8854 13163 -8842 se
rect 6756 -8917 6762 -8865
rect 6814 -8897 6829 -8865
rect 6881 -8897 6896 -8865
rect 6948 -8897 6963 -8865
rect 7015 -8897 7030 -8865
rect 7082 -8897 7096 -8865
rect 6822 -8917 6829 -8897
rect 7082 -8917 7088 -8897
rect 7148 -8917 7154 -8865
rect 6756 -8933 6766 -8917
rect 6822 -8933 6847 -8917
rect 6903 -8933 6928 -8917
rect 6984 -8933 7008 -8917
rect 7064 -8933 7088 -8917
rect 7144 -8933 7154 -8917
rect 6756 -8985 6762 -8933
rect 6822 -8953 6829 -8933
rect 7082 -8953 7088 -8933
rect 6814 -8985 6829 -8953
rect 6881 -8985 6896 -8953
rect 6948 -8985 6963 -8953
rect 7015 -8985 7030 -8953
rect 7082 -8985 7096 -8953
rect 7148 -8985 7154 -8933
<< rmetal2 >>
rect 2961 5312 2963 5364
<< via2 >>
rect 804 15831 856 15880
rect 856 15831 860 15880
rect 804 15824 860 15831
rect 884 15831 888 15880
rect 888 15831 940 15880
rect 884 15824 940 15831
rect 964 15831 972 15880
rect 972 15831 1020 15880
rect 964 15824 1020 15831
rect 804 15752 856 15793
rect 856 15752 860 15793
rect 804 15737 860 15752
rect 884 15752 888 15793
rect 888 15752 940 15793
rect 884 15737 940 15752
rect 964 15752 972 15793
rect 972 15752 1020 15793
rect 964 15737 1020 15752
rect 804 15673 856 15706
rect 856 15673 860 15706
rect 804 15650 860 15673
rect 884 15673 888 15706
rect 888 15673 940 15706
rect 884 15650 940 15673
rect 964 15673 972 15706
rect 972 15673 1020 15706
rect 964 15650 1020 15673
rect 804 15594 856 15618
rect 856 15594 860 15618
rect 804 15562 860 15594
rect 884 15594 888 15618
rect 888 15594 940 15618
rect 884 15562 940 15594
rect 964 15594 972 15618
rect 972 15594 1020 15618
rect 964 15562 1020 15594
rect 22995 7122 23051 7149
rect 22995 7093 23013 7122
rect 23013 7093 23051 7122
rect 22995 7058 23051 7069
rect 22995 7013 23013 7058
rect 23013 7013 23051 7058
rect 6343 6480 6391 6529
rect 6391 6480 6399 6529
rect 6425 6480 6457 6529
rect 6457 6480 6471 6529
rect 6471 6480 6481 6529
rect 6507 6480 6523 6529
rect 6523 6480 6537 6529
rect 6537 6480 6563 6529
rect 6589 6480 6603 6529
rect 6603 6480 6645 6529
rect 6671 6480 6720 6529
rect 6720 6480 6727 6529
rect 6753 6480 6785 6529
rect 6785 6480 6798 6529
rect 6798 6480 6809 6529
rect 6835 6480 6850 6529
rect 6850 6480 6863 6529
rect 6863 6480 6891 6529
rect 6917 6480 6928 6529
rect 6928 6480 6973 6529
rect 6999 6480 7045 6529
rect 7045 6480 7055 6529
rect 7081 6480 7110 6529
rect 7110 6480 7123 6529
rect 7123 6480 7137 6529
rect 7163 6480 7175 6529
rect 7175 6480 7188 6529
rect 7188 6480 7219 6529
rect 7245 6480 7253 6529
rect 7253 6480 7301 6529
rect 7326 6480 7370 6529
rect 7370 6480 7382 6529
rect 7407 6480 7435 6529
rect 7435 6480 7448 6529
rect 7448 6480 7463 6529
rect 7488 6480 7500 6529
rect 7500 6480 7513 6529
rect 7513 6480 7544 6529
rect 7569 6480 7578 6529
rect 7578 6480 7625 6529
rect 6343 6473 6399 6480
rect 6425 6473 6481 6480
rect 6507 6473 6563 6480
rect 6589 6473 6645 6480
rect 6671 6473 6727 6480
rect 6753 6473 6809 6480
rect 6835 6473 6891 6480
rect 6917 6473 6973 6480
rect 6999 6473 7055 6480
rect 7081 6473 7137 6480
rect 7163 6473 7219 6480
rect 7245 6473 7301 6480
rect 7326 6473 7382 6480
rect 7407 6473 7463 6480
rect 7488 6473 7544 6480
rect 7569 6473 7625 6480
rect 6343 6416 6399 6421
rect 6425 6416 6481 6421
rect 6507 6416 6563 6421
rect 6589 6416 6645 6421
rect 6671 6416 6727 6421
rect 6753 6416 6809 6421
rect 6835 6416 6891 6421
rect 6917 6416 6973 6421
rect 6999 6416 7055 6421
rect 7081 6416 7137 6421
rect 7163 6416 7219 6421
rect 7245 6416 7301 6421
rect 7326 6416 7382 6421
rect 7407 6416 7463 6421
rect 7488 6416 7544 6421
rect 7569 6416 7625 6421
rect 6343 6365 6391 6416
rect 6391 6365 6399 6416
rect 6425 6365 6457 6416
rect 6457 6365 6471 6416
rect 6471 6365 6481 6416
rect 6507 6365 6523 6416
rect 6523 6365 6537 6416
rect 6537 6365 6563 6416
rect 6589 6365 6603 6416
rect 6603 6365 6645 6416
rect 6671 6365 6720 6416
rect 6720 6365 6727 6416
rect 6753 6365 6785 6416
rect 6785 6365 6798 6416
rect 6798 6365 6809 6416
rect 6835 6365 6850 6416
rect 6850 6365 6863 6416
rect 6863 6365 6891 6416
rect 6917 6365 6928 6416
rect 6928 6365 6973 6416
rect 6999 6365 7045 6416
rect 7045 6365 7055 6416
rect 7081 6365 7110 6416
rect 7110 6365 7123 6416
rect 7123 6365 7137 6416
rect 7163 6365 7175 6416
rect 7175 6365 7188 6416
rect 7188 6365 7219 6416
rect 7245 6365 7253 6416
rect 7253 6365 7301 6416
rect 7326 6365 7370 6416
rect 7370 6365 7382 6416
rect 7407 6365 7435 6416
rect 7435 6365 7448 6416
rect 7448 6365 7463 6416
rect 7488 6365 7500 6416
rect 7500 6365 7513 6416
rect 7513 6365 7544 6416
rect 7569 6365 7578 6416
rect 7578 6365 7625 6416
rect 12521 6473 12577 6529
rect 12606 6473 12662 6529
rect 12691 6473 12747 6529
rect 12776 6473 12832 6529
rect 12860 6473 12916 6529
rect 12944 6473 13000 6529
rect 13028 6473 13084 6529
rect 12521 6365 12577 6421
rect 12606 6365 12662 6421
rect 12691 6365 12747 6421
rect 12776 6365 12832 6421
rect 12860 6365 12916 6421
rect 12944 6365 13000 6421
rect 13028 6365 13084 6421
rect 14328 6473 14384 6529
rect 14424 6473 14480 6529
rect 14519 6473 14575 6529
rect 14328 6365 14384 6421
rect 14424 6365 14480 6421
rect 14519 6365 14575 6421
rect 18363 6480 18411 6529
rect 18411 6480 18419 6529
rect 18444 6480 18480 6529
rect 18480 6480 18497 6529
rect 18497 6480 18500 6529
rect 18525 6480 18549 6529
rect 18549 6480 18565 6529
rect 18565 6480 18581 6529
rect 18606 6480 18617 6529
rect 18617 6480 18633 6529
rect 18633 6480 18662 6529
rect 18687 6480 18701 6529
rect 18701 6480 18743 6529
rect 18768 6480 18769 6529
rect 18769 6480 18821 6529
rect 18821 6480 18824 6529
rect 18849 6480 18889 6529
rect 18889 6480 18905 6529
rect 18929 6480 18957 6529
rect 18957 6480 18973 6529
rect 18973 6480 18985 6529
rect 19009 6480 19025 6529
rect 19025 6480 19041 6529
rect 19041 6480 19065 6529
rect 19089 6480 19093 6529
rect 19093 6480 19109 6529
rect 19109 6480 19145 6529
rect 19169 6480 19177 6529
rect 19177 6480 19225 6529
rect 18363 6473 18419 6480
rect 18444 6473 18500 6480
rect 18525 6473 18581 6480
rect 18606 6473 18662 6480
rect 18687 6473 18743 6480
rect 18768 6473 18824 6480
rect 18849 6473 18905 6480
rect 18929 6473 18985 6480
rect 19009 6473 19065 6480
rect 19089 6473 19145 6480
rect 19169 6473 19225 6480
rect 18363 6416 18419 6421
rect 18444 6416 18500 6421
rect 18525 6416 18581 6421
rect 18606 6416 18662 6421
rect 18687 6416 18743 6421
rect 18768 6416 18824 6421
rect 18849 6416 18905 6421
rect 18929 6416 18985 6421
rect 19009 6416 19065 6421
rect 19089 6416 19145 6421
rect 19169 6416 19225 6421
rect 18363 6365 18411 6416
rect 18411 6365 18419 6416
rect 18444 6365 18480 6416
rect 18480 6365 18497 6416
rect 18497 6365 18500 6416
rect 18525 6365 18549 6416
rect 18549 6365 18565 6416
rect 18565 6365 18581 6416
rect 18606 6365 18617 6416
rect 18617 6365 18633 6416
rect 18633 6365 18662 6416
rect 18687 6365 18701 6416
rect 18701 6365 18743 6416
rect 18768 6365 18769 6416
rect 18769 6365 18821 6416
rect 18821 6365 18824 6416
rect 18849 6365 18889 6416
rect 18889 6365 18905 6416
rect 18929 6365 18957 6416
rect 18957 6365 18973 6416
rect 18973 6365 18985 6416
rect 19009 6365 19025 6416
rect 19025 6365 19041 6416
rect 19041 6365 19065 6416
rect 19089 6365 19093 6416
rect 19093 6365 19109 6416
rect 19109 6365 19145 6416
rect 19169 6365 19177 6416
rect 19177 6365 19225 6416
rect 20202 6480 20250 6529
rect 20250 6480 20258 6529
rect 20283 6480 20319 6529
rect 20319 6480 20336 6529
rect 20336 6480 20339 6529
rect 20364 6480 20388 6529
rect 20388 6480 20404 6529
rect 20404 6480 20420 6529
rect 20445 6480 20456 6529
rect 20456 6480 20472 6529
rect 20472 6480 20501 6529
rect 20526 6480 20540 6529
rect 20540 6480 20582 6529
rect 20607 6480 20608 6529
rect 20608 6480 20660 6529
rect 20660 6480 20663 6529
rect 20688 6480 20728 6529
rect 20728 6480 20744 6529
rect 20768 6480 20796 6529
rect 20796 6480 20812 6529
rect 20812 6480 20824 6529
rect 20848 6480 20864 6529
rect 20864 6480 20880 6529
rect 20880 6480 20904 6529
rect 20928 6480 20932 6529
rect 20932 6480 20948 6529
rect 20948 6480 20984 6529
rect 21008 6480 21016 6529
rect 21016 6480 21064 6529
rect 20202 6473 20258 6480
rect 20283 6473 20339 6480
rect 20364 6473 20420 6480
rect 20445 6473 20501 6480
rect 20526 6473 20582 6480
rect 20607 6473 20663 6480
rect 20688 6473 20744 6480
rect 20768 6473 20824 6480
rect 20848 6473 20904 6480
rect 20928 6473 20984 6480
rect 21008 6473 21064 6480
rect 20202 6416 20258 6421
rect 20283 6416 20339 6421
rect 20364 6416 20420 6421
rect 20445 6416 20501 6421
rect 20526 6416 20582 6421
rect 20607 6416 20663 6421
rect 20688 6416 20744 6421
rect 20768 6416 20824 6421
rect 20848 6416 20904 6421
rect 20928 6416 20984 6421
rect 21008 6416 21064 6421
rect 20202 6365 20250 6416
rect 20250 6365 20258 6416
rect 20283 6365 20319 6416
rect 20319 6365 20336 6416
rect 20336 6365 20339 6416
rect 20364 6365 20388 6416
rect 20388 6365 20404 6416
rect 20404 6365 20420 6416
rect 20445 6365 20456 6416
rect 20456 6365 20472 6416
rect 20472 6365 20501 6416
rect 20526 6365 20540 6416
rect 20540 6365 20582 6416
rect 20607 6365 20608 6416
rect 20608 6365 20660 6416
rect 20660 6365 20663 6416
rect 20688 6365 20728 6416
rect 20728 6365 20744 6416
rect 20768 6365 20796 6416
rect 20796 6365 20812 6416
rect 20812 6365 20824 6416
rect 20848 6365 20864 6416
rect 20864 6365 20880 6416
rect 20880 6365 20904 6416
rect 20928 6365 20932 6416
rect 20932 6365 20948 6416
rect 20948 6365 20984 6416
rect 21008 6365 21016 6416
rect 21016 6365 21064 6416
rect 22985 6480 23033 6529
rect 23033 6480 23041 6529
rect 22985 6473 23041 6480
rect 23065 6480 23072 6529
rect 23072 6480 23121 6529
rect 23065 6473 23121 6480
rect 22985 6416 23041 6421
rect 22985 6365 23033 6416
rect 23033 6365 23041 6416
rect 23065 6416 23121 6421
rect 23065 6365 23072 6416
rect 23072 6365 23121 6416
rect 13720 -1459 13776 -1403
rect 13801 -1459 13857 -1403
rect 13882 -1459 13938 -1403
rect 13963 -1459 14019 -1403
rect 14044 -1459 14100 -1403
rect 14125 -1459 14181 -1403
rect 14206 -1459 14262 -1403
rect 14286 -1459 14342 -1403
rect 14366 -1459 14422 -1403
rect 14446 -1459 14502 -1403
rect 14526 -1459 14582 -1403
rect 18358 -1409 18414 -1353
rect 18439 -1409 18495 -1353
rect 18520 -1409 18576 -1353
rect 18601 -1409 18657 -1353
rect 18682 -1409 18738 -1353
rect 18763 -1409 18819 -1353
rect 18844 -1409 18900 -1353
rect 18924 -1409 18980 -1353
rect 19004 -1409 19060 -1353
rect 19084 -1409 19140 -1353
rect 19164 -1409 19220 -1353
rect 18358 -1470 18414 -1461
rect 18439 -1470 18495 -1461
rect 18520 -1470 18576 -1461
rect 18601 -1470 18657 -1461
rect 18682 -1470 18738 -1461
rect 18763 -1470 18819 -1461
rect 18844 -1470 18900 -1461
rect 18924 -1470 18980 -1461
rect 19004 -1470 19060 -1461
rect 19084 -1470 19140 -1461
rect 19164 -1470 19220 -1461
rect 18358 -1517 18407 -1470
rect 18407 -1517 18414 -1470
rect 18439 -1517 18475 -1470
rect 18475 -1517 18491 -1470
rect 18491 -1517 18495 -1470
rect 18520 -1517 18543 -1470
rect 18543 -1517 18559 -1470
rect 18559 -1517 18576 -1470
rect 18601 -1517 18611 -1470
rect 18611 -1517 18627 -1470
rect 18627 -1517 18657 -1470
rect 18682 -1517 18695 -1470
rect 18695 -1517 18738 -1470
rect 18763 -1517 18815 -1470
rect 18815 -1517 18819 -1470
rect 18844 -1517 18883 -1470
rect 18883 -1517 18899 -1470
rect 18899 -1517 18900 -1470
rect 18924 -1517 18951 -1470
rect 18951 -1517 18967 -1470
rect 18967 -1517 18980 -1470
rect 19004 -1517 19019 -1470
rect 19019 -1517 19035 -1470
rect 19035 -1517 19060 -1470
rect 19084 -1517 19087 -1470
rect 19087 -1517 19103 -1470
rect 19103 -1517 19140 -1470
rect 19164 -1517 19171 -1470
rect 19171 -1517 19220 -1470
rect 20199 -1409 20255 -1353
rect 20280 -1409 20336 -1353
rect 20361 -1409 20417 -1353
rect 20442 -1409 20498 -1353
rect 20523 -1409 20579 -1353
rect 20604 -1409 20660 -1353
rect 20685 -1409 20741 -1353
rect 20765 -1409 20821 -1353
rect 20845 -1409 20901 -1353
rect 20925 -1409 20981 -1353
rect 21005 -1409 21061 -1353
rect 20199 -1470 20255 -1461
rect 20280 -1470 20336 -1461
rect 20361 -1470 20417 -1461
rect 20442 -1470 20498 -1461
rect 20523 -1470 20579 -1461
rect 20604 -1470 20660 -1461
rect 20685 -1470 20741 -1461
rect 20765 -1470 20821 -1461
rect 20845 -1470 20901 -1461
rect 20925 -1470 20981 -1461
rect 21005 -1470 21061 -1461
rect 20199 -1517 20248 -1470
rect 20248 -1517 20255 -1470
rect 20280 -1517 20316 -1470
rect 20316 -1517 20332 -1470
rect 20332 -1517 20336 -1470
rect 20361 -1517 20384 -1470
rect 20384 -1517 20400 -1470
rect 20400 -1517 20417 -1470
rect 20442 -1517 20452 -1470
rect 20452 -1517 20468 -1470
rect 20468 -1517 20498 -1470
rect 20523 -1517 20536 -1470
rect 20536 -1517 20579 -1470
rect 20604 -1517 20656 -1470
rect 20656 -1517 20660 -1470
rect 20685 -1517 20724 -1470
rect 20724 -1517 20740 -1470
rect 20740 -1517 20741 -1470
rect 20765 -1517 20792 -1470
rect 20792 -1517 20808 -1470
rect 20808 -1517 20821 -1470
rect 20845 -1517 20860 -1470
rect 20860 -1517 20876 -1470
rect 20876 -1517 20901 -1470
rect 20925 -1517 20928 -1470
rect 20928 -1517 20944 -1470
rect 20944 -1517 20981 -1470
rect 21005 -1517 21012 -1470
rect 21012 -1517 21061 -1470
rect 6766 -7075 6814 -7056
rect 6814 -7075 6822 -7056
rect 6847 -7075 6881 -7056
rect 6881 -7075 6896 -7056
rect 6896 -7075 6903 -7056
rect 6928 -7075 6948 -7056
rect 6948 -7075 6963 -7056
rect 6963 -7075 6984 -7056
rect 7008 -7075 7015 -7056
rect 7015 -7075 7030 -7056
rect 7030 -7075 7064 -7056
rect 7088 -7075 7096 -7056
rect 7096 -7075 7144 -7056
rect 6766 -7091 6822 -7075
rect 6847 -7091 6903 -7075
rect 6928 -7091 6984 -7075
rect 7008 -7091 7064 -7075
rect 7088 -7091 7144 -7075
rect 6766 -7112 6814 -7091
rect 6814 -7112 6822 -7091
rect 6847 -7112 6881 -7091
rect 6881 -7112 6896 -7091
rect 6896 -7112 6903 -7091
rect 6928 -7112 6948 -7091
rect 6948 -7112 6963 -7091
rect 6963 -7112 6984 -7091
rect 7008 -7112 7015 -7091
rect 7015 -7112 7030 -7091
rect 7030 -7112 7064 -7091
rect 7088 -7112 7096 -7091
rect 7096 -7112 7144 -7091
rect 3167 -7396 3223 -7370
rect 3167 -7426 3216 -7396
rect 3216 -7426 3223 -7396
rect 3167 -7506 3223 -7450
rect 12645 -7401 12701 -7399
rect 12768 -7401 12824 -7399
rect 12891 -7401 12947 -7399
rect 13013 -7401 13069 -7399
rect 12645 -7453 12647 -7401
rect 12647 -7453 12699 -7401
rect 12699 -7453 12701 -7401
rect 12768 -7453 12791 -7401
rect 12791 -7453 12824 -7401
rect 12891 -7453 12922 -7401
rect 12922 -7453 12947 -7401
rect 13013 -7453 13065 -7401
rect 13065 -7453 13069 -7401
rect 12645 -7455 12701 -7453
rect 12768 -7455 12824 -7453
rect 12891 -7455 12947 -7453
rect 13013 -7455 13069 -7453
rect 12645 -7505 12701 -7503
rect 12768 -7505 12824 -7503
rect 12891 -7505 12947 -7503
rect 13013 -7505 13069 -7503
rect 12645 -7557 12647 -7505
rect 12647 -7557 12699 -7505
rect 12699 -7557 12701 -7505
rect 12768 -7557 12791 -7505
rect 12791 -7557 12824 -7505
rect 12891 -7557 12922 -7505
rect 12922 -7557 12947 -7505
rect 13013 -7557 13065 -7505
rect 13065 -7557 13069 -7505
rect 12645 -7559 12701 -7557
rect 12768 -7559 12824 -7557
rect 12891 -7559 12947 -7557
rect 13013 -7559 13069 -7557
rect 8274 -7615 8330 -7613
rect 8371 -7615 8427 -7613
rect 8467 -7615 8523 -7613
rect 8274 -7667 8285 -7615
rect 8285 -7667 8330 -7615
rect 8371 -7667 8377 -7615
rect 8377 -7667 8427 -7615
rect 8467 -7667 8469 -7615
rect 8469 -7667 8521 -7615
rect 8521 -7667 8523 -7615
rect 8274 -7669 8330 -7667
rect 8371 -7669 8427 -7667
rect 8467 -7669 8523 -7667
rect 12645 -7609 12701 -7607
rect 12768 -7609 12824 -7607
rect 12891 -7609 12947 -7607
rect 13013 -7609 13069 -7607
rect 12645 -7661 12647 -7609
rect 12647 -7661 12699 -7609
rect 12699 -7661 12701 -7609
rect 12768 -7661 12791 -7609
rect 12791 -7661 12824 -7609
rect 12891 -7661 12922 -7609
rect 12922 -7661 12947 -7609
rect 13013 -7661 13065 -7609
rect 13065 -7661 13069 -7609
rect 12645 -7663 12701 -7661
rect 12768 -7663 12824 -7661
rect 12891 -7663 12947 -7661
rect 13013 -7663 13069 -7661
rect 5141 -8285 5197 -8270
rect 5252 -8285 5308 -8270
rect 5363 -8285 5419 -8270
rect 5141 -8326 5151 -8285
rect 5151 -8326 5197 -8285
rect 5252 -8326 5302 -8285
rect 5302 -8326 5308 -8285
rect 5363 -8326 5400 -8285
rect 5400 -8326 5419 -8285
rect 5141 -8359 5197 -8354
rect 5252 -8359 5308 -8354
rect 5363 -8359 5419 -8354
rect 5141 -8410 5151 -8359
rect 5151 -8410 5197 -8359
rect 5252 -8410 5302 -8359
rect 5302 -8410 5308 -8359
rect 5363 -8410 5400 -8359
rect 5400 -8410 5419 -8359
rect 5141 -8485 5151 -8438
rect 5151 -8485 5197 -8438
rect 5252 -8485 5302 -8438
rect 5302 -8485 5308 -8438
rect 5363 -8485 5400 -8438
rect 5400 -8485 5419 -8438
rect 5141 -8494 5197 -8485
rect 5252 -8494 5308 -8485
rect 5363 -8494 5419 -8485
rect 5593 -8339 5597 -8287
rect 5597 -8339 5649 -8287
rect 5593 -8343 5649 -8339
rect 5681 -8343 5737 -8287
rect 5769 -8343 5825 -8287
rect 5856 -8343 5906 -8287
rect 5906 -8343 5912 -8287
rect 8374 -8355 8430 -8299
rect 5593 -8415 5649 -8411
rect 5593 -8467 5597 -8415
rect 5597 -8467 5649 -8415
rect 5681 -8467 5737 -8411
rect 5769 -8467 5825 -8411
rect 5856 -8467 5906 -8411
rect 5906 -8467 5912 -8411
rect 8374 -8435 8430 -8379
rect 6766 -8917 6814 -8897
rect 6814 -8917 6822 -8897
rect 6847 -8917 6881 -8897
rect 6881 -8917 6896 -8897
rect 6896 -8917 6903 -8897
rect 6928 -8917 6948 -8897
rect 6948 -8917 6963 -8897
rect 6963 -8917 6984 -8897
rect 7008 -8917 7015 -8897
rect 7015 -8917 7030 -8897
rect 7030 -8917 7064 -8897
rect 7088 -8917 7096 -8897
rect 7096 -8917 7144 -8897
rect 6766 -8933 6822 -8917
rect 6847 -8933 6903 -8917
rect 6928 -8933 6984 -8917
rect 7008 -8933 7064 -8917
rect 7088 -8933 7144 -8917
rect 6766 -8953 6814 -8933
rect 6814 -8953 6822 -8933
rect 6847 -8953 6881 -8933
rect 6881 -8953 6896 -8933
rect 6896 -8953 6903 -8933
rect 6928 -8953 6948 -8933
rect 6948 -8953 6963 -8933
rect 6963 -8953 6984 -8933
rect 7008 -8953 7015 -8933
rect 7015 -8953 7030 -8933
rect 7030 -8953 7064 -8933
rect 7088 -8953 7096 -8933
rect 7096 -8953 7144 -8933
<< metal3 >>
rect 707 15880 1309 16143
rect 707 15824 804 15880
rect 860 15824 884 15880
rect 940 15824 964 15880
rect 1020 15824 1309 15880
rect 707 15793 1309 15824
rect 707 15737 804 15793
rect 860 15737 884 15793
rect 940 15737 964 15793
rect 1020 15737 1309 15793
rect 707 15706 1309 15737
rect 707 15650 804 15706
rect 860 15650 884 15706
rect 940 15650 964 15706
rect 1020 15650 1309 15706
rect 707 15618 1309 15650
rect 707 15562 804 15618
rect 860 15562 884 15618
rect 940 15562 964 15618
rect 1020 15562 1309 15618
rect 707 -5992 1309 15562
rect 22980 7149 23126 7155
rect 22980 7093 22995 7149
rect 23051 7093 23126 7149
rect 22980 7069 23126 7093
rect 22980 7013 22995 7069
rect 23051 7013 23126 7069
rect 6333 6529 7703 6536
rect 6333 6473 6343 6529
rect 6399 6473 6425 6529
rect 6481 6473 6507 6529
rect 6563 6473 6589 6529
rect 6645 6473 6671 6529
rect 6727 6473 6753 6529
rect 6809 6473 6835 6529
rect 6891 6473 6917 6529
rect 6973 6473 6999 6529
rect 7055 6473 7081 6529
rect 7137 6473 7163 6529
rect 7219 6473 7245 6529
rect 7301 6473 7326 6529
rect 7382 6473 7407 6529
rect 7463 6473 7488 6529
rect 7544 6473 7569 6529
rect 7625 6473 7703 6529
rect 6333 6421 7703 6473
rect 6333 6365 6343 6421
rect 6399 6365 6425 6421
rect 6481 6365 6507 6421
rect 6563 6365 6589 6421
rect 6645 6365 6671 6421
rect 6727 6365 6753 6421
rect 6809 6365 6835 6421
rect 6891 6365 6917 6421
rect 6973 6365 6999 6421
rect 7055 6365 7081 6421
rect 7137 6365 7163 6421
rect 7219 6365 7245 6421
rect 7301 6365 7326 6421
rect 7382 6365 7407 6421
rect 7463 6365 7488 6421
rect 7544 6365 7569 6421
rect 7625 6365 7703 6421
rect 4343 -1244 5225 6257
rect 6333 5110 7703 6365
rect 12516 6529 13099 6536
rect 12516 6473 12521 6529
rect 12577 6473 12606 6529
rect 12662 6473 12691 6529
rect 12747 6473 12776 6529
rect 12832 6473 12860 6529
rect 12916 6473 12944 6529
rect 13000 6473 13028 6529
rect 13084 6473 13099 6529
rect 12516 6421 13099 6473
rect 12516 6365 12521 6421
rect 12577 6365 12606 6421
rect 12662 6365 12691 6421
rect 12747 6365 12776 6421
rect 12832 6365 12860 6421
rect 12916 6365 12944 6421
rect 13000 6365 13028 6421
rect 13084 6365 13099 6421
tri 12370 5517 12516 5663 se
rect 12516 5517 13099 6365
rect 14318 6529 14594 6536
rect 14318 6473 14328 6529
rect 14384 6473 14424 6529
rect 14480 6473 14519 6529
rect 14575 6473 14594 6529
rect 14318 6421 14594 6473
rect 14318 6365 14328 6421
rect 14384 6365 14424 6421
rect 14480 6365 14519 6421
rect 14575 6365 14594 6421
tri 7703 5110 8110 5517 sw
tri 12089 5236 12370 5517 se
rect 12370 5236 13099 5517
rect 6333 4949 8110 5110
tri 6333 4061 7221 4949 ne
rect 5985 -1788 6911 3088
rect 7221 -1244 8110 4949
tri 7345 -1353 7454 -1244 ne
rect 7454 -1353 8110 -1244
tri 11864 5011 12089 5236 se
rect 12089 5011 12753 5236
rect 11864 -1347 12753 5011
tri 12753 4890 13099 5236 nw
tri 13705 5010 14318 5623 se
rect 14318 5010 14594 6365
tri 11864 -1353 11870 -1347 ne
rect 11870 -1353 12753 -1347
tri 7454 -1362 7463 -1353 ne
rect 7463 -1578 8110 -1353
tri 11870 -1403 11920 -1353 ne
rect 11920 -1403 12753 -1353
tri 11920 -1418 11935 -1403 ne
rect 707 -6056 732 -5992
rect 796 -6056 812 -5992
rect 876 -6056 892 -5992
rect 956 -6056 972 -5992
rect 1036 -6056 1052 -5992
rect 1116 -6056 1132 -5992
rect 1196 -6056 1212 -5992
rect 1276 -6056 1309 -5992
rect 707 -6077 1309 -6056
rect 707 -6141 732 -6077
rect 796 -6141 812 -6077
rect 876 -6141 892 -6077
rect 956 -6141 972 -6077
rect 1036 -6141 1052 -6077
rect 1116 -6141 1132 -6077
rect 1196 -6141 1212 -6077
rect 1276 -6141 1309 -6077
rect 707 -6162 1309 -6141
rect 707 -6226 732 -6162
rect 796 -6226 812 -6162
rect 876 -6226 892 -6162
rect 956 -6226 972 -6162
rect 1036 -6226 1052 -6162
rect 1116 -6226 1132 -6162
rect 1196 -6226 1212 -6162
rect 1276 -6226 1309 -6162
rect 707 -6247 1309 -6226
rect 707 -6311 732 -6247
rect 796 -6311 812 -6247
rect 876 -6311 892 -6247
rect 956 -6311 972 -6247
rect 1036 -6311 1052 -6247
rect 1116 -6311 1132 -6247
rect 1196 -6311 1212 -6247
rect 1276 -6311 1309 -6247
rect 707 -6332 1309 -6311
rect 707 -6396 732 -6332
rect 796 -6396 812 -6332
rect 876 -6396 892 -6332
rect 956 -6396 972 -6332
rect 1036 -6396 1052 -6332
rect 1116 -6396 1132 -6332
rect 1196 -6396 1212 -6332
rect 1276 -6396 1309 -6332
rect 707 -6417 1309 -6396
rect 707 -6481 732 -6417
rect 796 -6481 812 -6417
rect 876 -6481 892 -6417
rect 956 -6481 972 -6417
rect 1036 -6481 1052 -6417
rect 1116 -6481 1132 -6417
rect 1196 -6481 1212 -6417
rect 1276 -6481 1309 -6417
rect 707 -6502 1309 -6481
rect 707 -6566 732 -6502
rect 796 -6566 812 -6502
rect 876 -6566 892 -6502
rect 956 -6566 972 -6502
rect 1036 -6566 1052 -6502
rect 1116 -6566 1132 -6502
rect 1196 -6566 1212 -6502
rect 1276 -6566 1309 -6502
rect 707 -6587 1309 -6566
rect 707 -6651 732 -6587
rect 796 -6651 812 -6587
rect 876 -6651 892 -6587
rect 956 -6651 972 -6587
rect 1036 -6651 1052 -6587
rect 1116 -6651 1132 -6587
rect 1196 -6651 1212 -6587
rect 1276 -6651 1309 -6587
rect 707 -6672 1309 -6651
rect 707 -6736 732 -6672
rect 796 -6736 812 -6672
rect 876 -6736 892 -6672
rect 956 -6736 972 -6672
rect 1036 -6736 1052 -6672
rect 1116 -6736 1132 -6672
rect 1196 -6736 1212 -6672
rect 1276 -6736 1309 -6672
rect 707 -6758 1309 -6736
rect 707 -6822 732 -6758
rect 796 -6822 812 -6758
rect 876 -6822 892 -6758
rect 956 -6822 972 -6758
rect 1036 -6822 1052 -6758
rect 1116 -6822 1132 -6758
rect 1196 -6822 1212 -6758
rect 1276 -6822 1309 -6758
rect 707 -6844 1309 -6822
rect 707 -6908 732 -6844
rect 796 -6908 812 -6844
rect 876 -6908 892 -6844
rect 956 -6908 972 -6844
rect 1036 -6908 1052 -6844
rect 1116 -6908 1132 -6844
rect 1196 -6908 1212 -6844
rect 1276 -6908 1309 -6844
rect 707 -6915 1309 -6908
rect 3154 -7370 3240 -1868
rect 11935 -2429 12753 -1403
rect 13705 -1403 14594 5010
rect 13705 -1459 13720 -1403
rect 13776 -1459 13801 -1403
rect 13857 -1459 13882 -1403
rect 13938 -1459 13963 -1403
rect 14019 -1459 14044 -1403
rect 14100 -1459 14125 -1403
rect 14181 -1459 14206 -1403
rect 14262 -1459 14286 -1403
rect 14342 -1459 14366 -1403
rect 14422 -1459 14446 -1403
rect 14502 -1459 14526 -1403
rect 14582 -1459 14594 -1403
rect 13705 -1464 14594 -1459
rect 18348 6529 19237 6536
rect 18348 6473 18363 6529
rect 18419 6473 18444 6529
rect 18500 6473 18525 6529
rect 18581 6473 18606 6529
rect 18662 6473 18687 6529
rect 18743 6473 18768 6529
rect 18824 6473 18849 6529
rect 18905 6473 18929 6529
rect 18985 6473 19009 6529
rect 19065 6473 19089 6529
rect 19145 6473 19169 6529
rect 19225 6473 19237 6529
rect 18348 6421 19237 6473
rect 18348 6365 18363 6421
rect 18419 6365 18444 6421
rect 18500 6365 18525 6421
rect 18581 6365 18606 6421
rect 18662 6365 18687 6421
rect 18743 6365 18768 6421
rect 18824 6365 18849 6421
rect 18905 6365 18929 6421
rect 18985 6365 19009 6421
rect 19065 6365 19089 6421
rect 19145 6365 19169 6421
rect 19225 6365 19237 6421
rect 18348 -1353 19237 6365
rect 18348 -1409 18358 -1353
rect 18414 -1409 18439 -1353
rect 18495 -1409 18520 -1353
rect 18576 -1409 18601 -1353
rect 18657 -1409 18682 -1353
rect 18738 -1409 18763 -1353
rect 18819 -1409 18844 -1353
rect 18900 -1409 18924 -1353
rect 18980 -1409 19004 -1353
rect 19060 -1409 19084 -1353
rect 19140 -1409 19164 -1353
rect 19220 -1409 19237 -1353
rect 18348 -1461 19237 -1409
rect 18348 -1517 18358 -1461
rect 18414 -1517 18439 -1461
rect 18495 -1517 18520 -1461
rect 18576 -1517 18601 -1461
rect 18657 -1517 18682 -1461
rect 18738 -1517 18763 -1461
rect 18819 -1517 18844 -1461
rect 18900 -1517 18924 -1461
rect 18980 -1517 19004 -1461
rect 19060 -1517 19084 -1461
rect 19140 -1517 19164 -1461
rect 19220 -1517 19237 -1461
rect 18348 -1792 19237 -1517
rect 20189 6529 21078 6536
rect 20189 6473 20202 6529
rect 20258 6473 20283 6529
rect 20339 6473 20364 6529
rect 20420 6473 20445 6529
rect 20501 6473 20526 6529
rect 20582 6473 20607 6529
rect 20663 6473 20688 6529
rect 20744 6473 20768 6529
rect 20824 6473 20848 6529
rect 20904 6473 20928 6529
rect 20984 6473 21008 6529
rect 21064 6473 21078 6529
rect 20189 6421 21078 6473
rect 20189 6365 20202 6421
rect 20258 6365 20283 6421
rect 20339 6365 20364 6421
rect 20420 6365 20445 6421
rect 20501 6365 20526 6421
rect 20582 6365 20607 6421
rect 20663 6365 20688 6421
rect 20744 6365 20768 6421
rect 20824 6365 20848 6421
rect 20904 6365 20928 6421
rect 20984 6365 21008 6421
rect 21064 6365 21078 6421
rect 20189 -1353 21078 6365
rect 22980 6529 23126 7013
rect 22980 6473 22985 6529
rect 23041 6473 23065 6529
rect 23121 6473 23126 6529
rect 22980 6421 23126 6473
rect 22980 6365 22985 6421
rect 23041 6365 23065 6421
rect 23121 6365 23126 6421
rect 22980 1312 23126 6365
rect 20189 -1409 20199 -1353
rect 20255 -1409 20280 -1353
rect 20336 -1409 20361 -1353
rect 20417 -1409 20442 -1353
rect 20498 -1409 20523 -1353
rect 20579 -1409 20604 -1353
rect 20660 -1409 20685 -1353
rect 20741 -1409 20765 -1353
rect 20821 -1409 20845 -1353
rect 20901 -1409 20925 -1353
rect 20981 -1409 21005 -1353
rect 21061 -1409 21078 -1353
rect 20189 -1461 21078 -1409
rect 20189 -1517 20199 -1461
rect 20255 -1517 20280 -1461
rect 20336 -1517 20361 -1461
rect 20417 -1517 20442 -1461
rect 20498 -1517 20523 -1461
rect 20579 -1517 20604 -1461
rect 20660 -1517 20685 -1461
rect 20741 -1517 20765 -1461
rect 20821 -1517 20845 -1461
rect 20901 -1517 20925 -1461
rect 20981 -1517 21005 -1461
rect 21061 -1517 21078 -1461
rect 20189 -1795 21078 -1517
tri 11935 -2711 12217 -2429 ne
rect 12217 -2711 12753 -2429
tri 12753 -2711 13089 -2375 sw
tri 12217 -3126 12632 -2711 ne
rect 3154 -7426 3167 -7370
rect 3223 -7426 3240 -7370
rect 3154 -7450 3240 -7426
rect 3154 -7506 3167 -7450
rect 3223 -7506 3240 -7450
rect 3154 -7563 3240 -7506
rect 5068 -7455 5397 -7001
rect 6761 -7056 7149 -7021
rect 6761 -7112 6766 -7056
rect 6822 -7112 6847 -7056
rect 6903 -7112 6928 -7056
rect 6984 -7112 7008 -7056
rect 7064 -7112 7088 -7056
rect 7144 -7112 7149 -7056
tri 5397 -7455 5400 -7452 sw
rect 5068 -7503 5400 -7455
tri 5400 -7503 5448 -7455 sw
rect 5068 -7508 5448 -7503
tri 5448 -7508 5453 -7503 sw
rect 5068 -7559 5453 -7508
tri 5453 -7559 5504 -7508 sw
rect 5068 -7563 5504 -7559
tri 5504 -7563 5508 -7559 sw
rect 5068 -7587 5508 -7563
tri 5068 -7607 5088 -7587 ne
rect 5088 -7607 5508 -7587
tri 5508 -7607 5552 -7563 sw
tri 5088 -7613 5094 -7607 ne
rect 5094 -7613 5552 -7607
tri 5552 -7613 5558 -7607 sw
tri 5094 -7669 5150 -7613 ne
rect 5150 -7669 5558 -7613
tri 5558 -7669 5614 -7613 sw
tri 5150 -7972 5453 -7669 ne
rect 5453 -7972 5614 -7669
tri 5614 -7972 5917 -7669 sw
tri 5453 -8107 5588 -7972 ne
rect 5136 -8270 5424 -8265
rect 5136 -8326 5141 -8270
rect 5197 -8326 5252 -8270
rect 5308 -8326 5363 -8270
rect 5419 -8326 5424 -8270
rect 5136 -8354 5424 -8326
rect 5136 -8410 5141 -8354
rect 5197 -8410 5252 -8354
rect 5308 -8410 5363 -8354
rect 5419 -8410 5424 -8354
rect 5136 -8438 5424 -8410
rect 5136 -8494 5141 -8438
rect 5197 -8494 5252 -8438
rect 5308 -8494 5363 -8438
rect 5419 -8494 5424 -8438
rect 5588 -8287 5917 -7972
rect 5588 -8343 5593 -8287
rect 5649 -8343 5681 -8287
rect 5737 -8343 5769 -8287
rect 5825 -8343 5856 -8287
rect 5912 -8343 5917 -8287
rect 5588 -8411 5917 -8343
rect 5588 -8467 5593 -8411
rect 5649 -8467 5681 -8411
rect 5737 -8467 5769 -8411
rect 5825 -8467 5856 -8411
rect 5912 -8467 5917 -8411
rect 5588 -8472 5917 -8467
tri 6549 -8472 6581 -8440 se
rect 6581 -8472 6619 -8440
rect 5136 -8648 5424 -8494
tri 6425 -8596 6549 -8472 se
rect 6549 -8596 6619 -8472
tri 5424 -8648 5476 -8596 sw
tri 6373 -8648 6425 -8596 se
rect 6425 -8648 6619 -8596
rect 5136 -8714 6619 -8648
tri 5136 -8897 5319 -8714 ne
rect 5319 -8897 6619 -8714
tri 5319 -8936 5358 -8897 ne
rect 5358 -8936 6619 -8897
tri 6379 -8953 6396 -8936 ne
rect 6396 -8953 6619 -8936
tri 6396 -9138 6581 -8953 ne
rect 6581 -9138 6619 -8953
rect 6761 -8897 7149 -7112
rect 12632 -7399 13089 -2711
rect 12632 -7455 12645 -7399
rect 12701 -7455 12768 -7399
rect 12824 -7455 12891 -7399
rect 12947 -7455 13013 -7399
rect 13069 -7455 13089 -7399
rect 12632 -7503 13089 -7455
rect 12632 -7559 12645 -7503
rect 12701 -7559 12768 -7503
rect 12824 -7559 12891 -7503
rect 12947 -7559 13013 -7503
rect 13069 -7559 13089 -7503
rect 12632 -7607 13089 -7559
rect 8269 -7613 8528 -7608
rect 8269 -7669 8274 -7613
rect 8330 -7669 8371 -7613
rect 8427 -7669 8467 -7613
rect 8523 -7669 8528 -7613
rect 12632 -7663 12645 -7607
rect 12701 -7663 12768 -7607
rect 12824 -7663 12891 -7607
rect 12947 -7663 13013 -7607
rect 13069 -7663 13089 -7607
rect 12632 -7669 13089 -7663
rect 8269 -7689 8528 -7669
tri 8269 -7764 8344 -7689 ne
rect 8344 -8183 8460 -7689
tri 8460 -7757 8528 -7689 nw
rect 8344 -8299 8460 -8294
rect 8344 -8355 8374 -8299
rect 8430 -8355 8460 -8299
rect 8344 -8379 8460 -8355
rect 8344 -8435 8374 -8379
rect 8430 -8435 8460 -8379
rect 8344 -8440 8460 -8435
rect 6761 -8953 6766 -8897
rect 6822 -8953 6847 -8897
rect 6903 -8953 6928 -8897
rect 6984 -8953 7008 -8897
rect 7064 -8953 7088 -8897
rect 7144 -8953 7149 -8897
rect 6761 -8988 7149 -8953
<< via3 >>
rect 732 -6056 796 -5992
rect 812 -6056 876 -5992
rect 892 -6056 956 -5992
rect 972 -6056 1036 -5992
rect 1052 -6056 1116 -5992
rect 1132 -6056 1196 -5992
rect 1212 -6056 1276 -5992
rect 732 -6141 796 -6077
rect 812 -6141 876 -6077
rect 892 -6141 956 -6077
rect 972 -6141 1036 -6077
rect 1052 -6141 1116 -6077
rect 1132 -6141 1196 -6077
rect 1212 -6141 1276 -6077
rect 732 -6226 796 -6162
rect 812 -6226 876 -6162
rect 892 -6226 956 -6162
rect 972 -6226 1036 -6162
rect 1052 -6226 1116 -6162
rect 1132 -6226 1196 -6162
rect 1212 -6226 1276 -6162
rect 732 -6311 796 -6247
rect 812 -6311 876 -6247
rect 892 -6311 956 -6247
rect 972 -6311 1036 -6247
rect 1052 -6311 1116 -6247
rect 1132 -6311 1196 -6247
rect 1212 -6311 1276 -6247
rect 732 -6396 796 -6332
rect 812 -6396 876 -6332
rect 892 -6396 956 -6332
rect 972 -6396 1036 -6332
rect 1052 -6396 1116 -6332
rect 1132 -6396 1196 -6332
rect 1212 -6396 1276 -6332
rect 732 -6481 796 -6417
rect 812 -6481 876 -6417
rect 892 -6481 956 -6417
rect 972 -6481 1036 -6417
rect 1052 -6481 1116 -6417
rect 1132 -6481 1196 -6417
rect 1212 -6481 1276 -6417
rect 732 -6566 796 -6502
rect 812 -6566 876 -6502
rect 892 -6566 956 -6502
rect 972 -6566 1036 -6502
rect 1052 -6566 1116 -6502
rect 1132 -6566 1196 -6502
rect 1212 -6566 1276 -6502
rect 732 -6651 796 -6587
rect 812 -6651 876 -6587
rect 892 -6651 956 -6587
rect 972 -6651 1036 -6587
rect 1052 -6651 1116 -6587
rect 1132 -6651 1196 -6587
rect 1212 -6651 1276 -6587
rect 732 -6736 796 -6672
rect 812 -6736 876 -6672
rect 892 -6736 956 -6672
rect 972 -6736 1036 -6672
rect 1052 -6736 1116 -6672
rect 1132 -6736 1196 -6672
rect 1212 -6736 1276 -6672
rect 732 -6822 796 -6758
rect 812 -6822 876 -6758
rect 892 -6822 956 -6758
rect 972 -6822 1036 -6758
rect 1052 -6822 1116 -6758
rect 1132 -6822 1196 -6758
rect 1212 -6822 1276 -6758
rect 732 -6908 796 -6844
rect 812 -6908 876 -6844
rect 892 -6908 956 -6844
rect 972 -6908 1036 -6844
rect 1052 -6908 1116 -6844
rect 1132 -6908 1196 -6844
rect 1212 -6908 1276 -6844
<< metal4 >>
rect 731 -5992 1277 -5991
rect 731 -6056 732 -5992
rect 796 -6056 812 -5992
rect 876 -6056 892 -5992
rect 956 -6056 972 -5992
rect 1036 -6056 1052 -5992
rect 1116 -6056 1132 -5992
rect 1196 -6056 1212 -5992
rect 1276 -6056 1277 -5992
rect 731 -6077 1277 -6056
rect 731 -6141 732 -6077
rect 796 -6141 812 -6077
rect 876 -6141 892 -6077
rect 956 -6141 972 -6077
rect 1036 -6141 1052 -6077
rect 1116 -6141 1132 -6077
rect 1196 -6141 1212 -6077
rect 1276 -6141 1277 -6077
rect 731 -6162 1277 -6141
rect 731 -6226 732 -6162
rect 796 -6226 812 -6162
rect 876 -6226 892 -6162
rect 956 -6226 972 -6162
rect 1036 -6226 1052 -6162
rect 1116 -6226 1132 -6162
rect 1196 -6226 1212 -6162
rect 1276 -6226 1277 -6162
rect 731 -6247 1277 -6226
rect 731 -6311 732 -6247
rect 796 -6311 812 -6247
rect 876 -6311 892 -6247
rect 956 -6311 972 -6247
rect 1036 -6311 1052 -6247
rect 1116 -6311 1132 -6247
rect 1196 -6311 1212 -6247
rect 1276 -6311 1277 -6247
rect 731 -6332 1277 -6311
rect 731 -6396 732 -6332
rect 796 -6396 812 -6332
rect 876 -6396 892 -6332
rect 956 -6396 972 -6332
rect 1036 -6396 1052 -6332
rect 1116 -6396 1132 -6332
rect 1196 -6396 1212 -6332
rect 1276 -6396 1277 -6332
rect 731 -6417 1277 -6396
rect 731 -6481 732 -6417
rect 796 -6481 812 -6417
rect 876 -6481 892 -6417
rect 956 -6481 972 -6417
rect 1036 -6481 1052 -6417
rect 1116 -6481 1132 -6417
rect 1196 -6481 1212 -6417
rect 1276 -6481 1277 -6417
rect 731 -6502 1277 -6481
rect 731 -6566 732 -6502
rect 796 -6566 812 -6502
rect 876 -6566 892 -6502
rect 956 -6566 972 -6502
rect 1036 -6566 1052 -6502
rect 1116 -6566 1132 -6502
rect 1196 -6566 1212 -6502
rect 1276 -6566 1277 -6502
rect 731 -6587 1277 -6566
rect 731 -6651 732 -6587
rect 796 -6651 812 -6587
rect 876 -6651 892 -6587
rect 956 -6651 972 -6587
rect 1036 -6651 1052 -6587
rect 1116 -6651 1132 -6587
rect 1196 -6651 1212 -6587
rect 1276 -6651 1277 -6587
rect 731 -6672 1277 -6651
rect 731 -6736 732 -6672
rect 796 -6736 812 -6672
rect 876 -6736 892 -6672
rect 956 -6736 972 -6672
rect 1036 -6736 1052 -6672
rect 1116 -6736 1132 -6672
rect 1196 -6736 1212 -6672
rect 1276 -6736 1277 -6672
rect 731 -6758 1277 -6736
rect 731 -6822 732 -6758
rect 796 -6822 812 -6758
rect 876 -6822 892 -6758
rect 956 -6822 972 -6758
rect 1036 -6822 1052 -6758
rect 1116 -6822 1132 -6758
rect 1196 -6822 1212 -6758
rect 1276 -6822 1277 -6758
rect 731 -6844 1277 -6822
rect 731 -6908 732 -6844
rect 796 -6908 812 -6844
rect 876 -6908 892 -6844
rect 956 -6908 972 -6844
rect 1036 -6908 1052 -6844
rect 1116 -6908 1132 -6844
rect 1196 -6908 1212 -6844
rect 1276 -6908 1277 -6844
rect 731 -6909 1277 -6908
use sky130_fd_io__gpio_ovtv2_hotswap_bias  sky130_fd_io__gpio_ovtv2_hotswap_bias_0
timestamp 1683767628
transform 1 0 1604 0 1 -769
box -1236 -1179 25744 7485
use sky130_fd_io__gpio_ovtv2_hotswap_guardrings  sky130_fd_io__gpio_ovtv2_hotswap_guardrings_0
timestamp 1683767628
transform 1 0 368 0 1 -1948
box 0 0 26980 8664
use sky130_fd_io__gpio_ovtv2_hotswap_nonoverlap_leak_fix  sky130_fd_io__gpio_ovtv2_hotswap_nonoverlap_leak_fix_0
timestamp 1683767628
transform 0 1 -5775 -1 0 6515
box -11144 5775 6448 12812
use sky130_fd_io__gpio_ovtv2_hotswap_pghs_i2c_fix  sky130_fd_io__gpio_ovtv2_hotswap_pghs_i2c_fix_0
timestamp 1683767628
transform 1 0 -114 0 1 -9106
box 174 25 27462 15822
use sky130_fd_io__gpio_ovtv2_hotswap_pug  sky130_fd_io__gpio_ovtv2_hotswap_pug_0
array 0 5 3220 0 0 494
timestamp 1683767628
transform 1 0 6184 0 -1 5161
box 0 0 3318 507
use sky130_fd_io__gpio_ovtv2_hotswap_pug_ovtfix  sky130_fd_io__gpio_ovtv2_hotswap_pug_ovtfix_0
timestamp 1683767628
transform 1 0 2964 0 -1 5161
box 0 0 3318 507
use sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias  sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_0
timestamp 1683767628
transform 1 0 2995 0 1 1299
box -2627 -3247 24353 5417
use sky130_fd_pr__m1short__example_55959141808175  sky130_fd_pr__m1short__example_55959141808175_0
timestamp 1683767628
transform 0 -1 23734 1 0 2839
box 0 0 1 1
use sky130_fd_pr__m1short__example_55959141808175  sky130_fd_pr__m1short__example_55959141808175_1
timestamp 1683767628
transform 1 0 23792 0 1 2731
box 0 0 1 1
use sky130_fd_pr__m2short__example_55959141808176  sky130_fd_pr__m2short__example_55959141808176_0
timestamp 1683767628
transform -1 0 2986 0 -1 5364
box 0 0 1 1
use sky130_fd_pr__res_generic_po__example_5595914180838  sky130_fd_pr__res_generic_po__example_5595914180838_0
timestamp 1683767628
transform 1 0 23066 0 1 7026
box 15 17 2025 18
use sky130_fd_pr__res_generic_po__example_5595914180838  sky130_fd_pr__res_generic_po__example_5595914180838_1
timestamp 1683767628
transform -1 0 25115 0 1 7252
box 15 17 2025 18
<< labels >>
flabel comment s 25602 5414 25602 5414 0 FreeSans 200 0 0 0 VCC_IO_SOFT
flabel comment s 3962 4965 3962 4965 0 FreeSans 1200 0 0 0 4
flabel comment s 7873 4997 7873 4997 0 FreeSans 1200 0 0 0 6
flabel comment s 9765 4982 9765 4982 0 FreeSans 1200 0 0 0 5
flabel comment s 13270 4997 13270 4997 0 FreeSans 1200 0 0 0 3
flabel comment s 16233 4995 16233 4995 0 FreeSans 1200 0 0 0 2
flabel comment s 19298 5004 19298 5004 0 FreeSans 1200 0 0 0 1
flabel comment s 23168 4994 23168 4994 0 FreeSans 400 0 0 0 0
flabel comment s 7182 4965 7182 4965 0 FreeSans 1200 0 0 0 4
flabel comment s 11093 4997 11093 4997 0 FreeSans 1200 0 0 0 6
flabel comment s 12985 4982 12985 4982 0 FreeSans 1200 0 0 0 5
flabel comment s 16490 4997 16490 4997 0 FreeSans 1200 0 0 0 3
flabel comment s 19453 4995 19453 4995 0 FreeSans 1200 0 0 0 2
flabel comment s 22518 5004 22518 5004 0 FreeSans 1200 0 0 0 1
flabel comment s 26388 4994 26388 4994 0 FreeSans 400 0 0 0 0
flabel comment s 25529 5245 25529 5245 0 FreeSans 400 0 0 0 TIE_HI
flabel comment s 16233 4995 16233 4995 0 FreeSans 1200 0 0 0 2
flabel comment s 13270 4997 13270 4997 0 FreeSans 1200 0 0 0 3
flabel comment s 9765 4982 9765 4982 0 FreeSans 1200 0 0 0 5
flabel comment s 3962 4965 3962 4965 0 FreeSans 1200 0 0 0 4
flabel comment s 7873 4997 7873 4997 0 FreeSans 1200 0 0 0 6
flabel comment s 19298 5004 19298 5004 0 FreeSans 1200 0 0 0 1
flabel comment s 23168 4994 23168 4994 0 FreeSans 1000 0 0 0 0
flabel metal1 s 1599 -420 1830 -249 3 FreeSans 520 0 0 0 VPB_DRVR
port 1 nsew
flabel metal1 s 22920 4594 22955 4626 3 FreeSans 200 0 0 0 PUG_H[0]
port 2 nsew
flabel metal1 s 19577 4535 19614 4566 3 FreeSans 200 0 0 0 PUG_H[1]
port 3 nsew
flabel metal1 s 16314 5174 16352 5209 3 FreeSans 200 0 0 0 PUG_H[2]
port 4 nsew
flabel metal1 s 13516 4397 13554 4433 3 FreeSans 200 0 0 0 PUG_H[3]
port 5 nsew
flabel metal1 s 2772 4742 2808 4774 3 FreeSans 200 0 0 0 PUG_H[4]
port 6 nsew
flabel metal1 s 9489 4897 9521 4929 3 FreeSans 200 0 0 0 PUG_H[5]
port 7 nsew
flabel metal1 s 7905 4467 7940 4499 3 FreeSans 200 0 0 0 PUG_H[6]
port 8 nsew
flabel metal1 s 932 12912 1002 13195 3 FreeSans 520 0 0 0 VSSD
port 9 nsew
flabel metal1 s 2451 947 2491 993 3 FreeSans 200 0 0 0 P2G
port 10 nsew
flabel metal1 s 10695 -8146 10784 -8092 3 FreeSans 200 0 0 0 OE_HS_H
port 11 nsew
flabel metal1 s 10423 -8162 10487 -8124 3 FreeSans 200 0 0 0 FORCE_H[1]
port 12 nsew
flabel metal1 s 11829 -8226 11889 -8194 3 FreeSans 200 0 0 0 OD_H
port 13 nsew
flabel metal1 s 7639 -8357 7738 -8311 3 FreeSans 200 0 0 0 VPWR_KA
port 14 nsew
flabel metal1 s 1753 5468 1936 5552 3 FreeSans 200 0 0 0 PAD_ESD
port 15 nsew
flabel metal1 s 684 -1792 930 -1613 3 FreeSans 520 0 0 0 VDDIO
port 16 nsew
flabel metal2 s 2004 765 2031 792 0 FreeSans 200 90 0 0 NGHS_H
port 18 nsew
flabel metal2 s 2671 5231 2723 5271 3 FreeSans 200 0 0 0 PGHS_H
port 19 nsew
flabel metal2 s 25570 6819 25721 6864 3 FreeSans 200 0 0 0 VCC_IO_SOFT
port 20 nsew
flabel metal2 s 26647 -5487 26930 -5417 3 FreeSans 520 90 0 0 VSSD
port 9 nsew
flabel metal2 s 8386 3591 8803 3697 3 FreeSans 520 0 0 0 PAD
port 21 nsew
<< properties >>
string GDS_END 40431348
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 40342612
<< end >>
