magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect 173 1122 1076 1664
rect 173 963 1598 1122
rect 179 956 1598 963
rect 1114 413 1559 956
rect 24705 -1927 25239 -1226
<< pwell >>
rect 239 1984 1020 2070
rect 254 1769 994 1984
rect 1200 93 1478 308
rect 255 7 1552 93
rect 24745 -1121 25202 -929
<< mvnmos >>
rect 333 1795 453 1935
rect 619 1795 739 1935
rect 795 1795 915 1935
rect 1279 142 1399 282
rect 24824 -1095 24944 -955
rect 25000 -1095 25120 -955
<< mvpmos >>
rect 333 1397 453 1597
rect 619 1397 739 1597
rect 795 1397 915 1597
rect 333 1129 453 1329
rect 619 1129 739 1329
rect 795 1129 915 1329
rect 1279 748 1399 948
rect 1279 480 1399 680
rect 24824 -1493 24944 -1293
rect 25000 -1493 25120 -1293
rect 24824 -1761 24944 -1561
rect 25000 -1761 25120 -1561
<< mvndiff >>
rect 280 1909 333 1935
rect 280 1875 288 1909
rect 322 1875 333 1909
rect 280 1841 333 1875
rect 280 1807 288 1841
rect 322 1807 333 1841
rect 280 1795 333 1807
rect 453 1909 506 1935
rect 453 1875 464 1909
rect 498 1875 506 1909
rect 453 1841 506 1875
rect 453 1807 464 1841
rect 498 1807 506 1841
rect 453 1795 506 1807
rect 566 1909 619 1935
rect 566 1875 574 1909
rect 608 1875 619 1909
rect 566 1841 619 1875
rect 566 1807 574 1841
rect 608 1807 619 1841
rect 566 1795 619 1807
rect 739 1795 795 1935
rect 915 1909 968 1935
rect 915 1875 926 1909
rect 960 1875 968 1909
rect 915 1841 968 1875
rect 915 1807 926 1841
rect 960 1807 968 1841
rect 915 1795 968 1807
rect 1226 270 1279 282
rect 1226 236 1234 270
rect 1268 236 1279 270
rect 1226 202 1279 236
rect 1226 168 1234 202
rect 1268 168 1279 202
rect 1226 142 1279 168
rect 1399 270 1452 282
rect 1399 236 1410 270
rect 1444 236 1452 270
rect 1399 202 1452 236
rect 1399 168 1410 202
rect 1444 168 1452 202
rect 1399 142 1452 168
rect 24771 -981 24824 -955
rect 24771 -1015 24779 -981
rect 24813 -1015 24824 -981
rect 24771 -1049 24824 -1015
rect 24771 -1083 24779 -1049
rect 24813 -1083 24824 -1049
rect 24771 -1095 24824 -1083
rect 24944 -981 25000 -955
rect 24944 -1015 24955 -981
rect 24989 -1015 25000 -981
rect 24944 -1049 25000 -1015
rect 24944 -1083 24955 -1049
rect 24989 -1083 25000 -1049
rect 24944 -1095 25000 -1083
rect 25120 -981 25176 -955
rect 25120 -1015 25131 -981
rect 25165 -1015 25176 -981
rect 25120 -1049 25176 -1015
rect 25120 -1083 25131 -1049
rect 25165 -1083 25176 -1049
rect 25120 -1095 25176 -1083
<< mvpdiff >>
rect 280 1579 333 1597
rect 280 1545 288 1579
rect 322 1545 333 1579
rect 280 1511 333 1545
rect 280 1477 288 1511
rect 322 1477 333 1511
rect 280 1443 333 1477
rect 280 1409 288 1443
rect 322 1409 333 1443
rect 280 1397 333 1409
rect 453 1579 506 1597
rect 453 1545 464 1579
rect 498 1545 506 1579
rect 453 1511 506 1545
rect 453 1477 464 1511
rect 498 1477 506 1511
rect 453 1443 506 1477
rect 453 1409 464 1443
rect 498 1409 506 1443
rect 453 1397 506 1409
rect 566 1579 619 1597
rect 566 1545 574 1579
rect 608 1545 619 1579
rect 566 1511 619 1545
rect 566 1477 574 1511
rect 608 1477 619 1511
rect 566 1443 619 1477
rect 566 1409 574 1443
rect 608 1409 619 1443
rect 566 1397 619 1409
rect 739 1579 795 1597
rect 739 1545 750 1579
rect 784 1545 795 1579
rect 739 1511 795 1545
rect 739 1477 750 1511
rect 784 1477 795 1511
rect 739 1443 795 1477
rect 739 1409 750 1443
rect 784 1409 795 1443
rect 739 1397 795 1409
rect 915 1579 968 1597
rect 915 1545 926 1579
rect 960 1545 968 1579
rect 915 1511 968 1545
rect 915 1477 926 1511
rect 960 1477 968 1511
rect 915 1443 968 1477
rect 915 1409 926 1443
rect 960 1409 968 1443
rect 915 1397 968 1409
rect 280 1317 333 1329
rect 280 1283 288 1317
rect 322 1283 333 1317
rect 280 1249 333 1283
rect 280 1215 288 1249
rect 322 1215 333 1249
rect 280 1181 333 1215
rect 280 1147 288 1181
rect 322 1147 333 1181
rect 280 1129 333 1147
rect 453 1317 506 1329
rect 453 1283 464 1317
rect 498 1283 506 1317
rect 453 1249 506 1283
rect 453 1215 464 1249
rect 498 1215 506 1249
rect 453 1181 506 1215
rect 453 1147 464 1181
rect 498 1147 506 1181
rect 453 1129 506 1147
rect 566 1317 619 1329
rect 566 1283 574 1317
rect 608 1283 619 1317
rect 566 1249 619 1283
rect 566 1215 574 1249
rect 608 1215 619 1249
rect 566 1181 619 1215
rect 566 1147 574 1181
rect 608 1147 619 1181
rect 566 1129 619 1147
rect 739 1317 795 1329
rect 739 1283 750 1317
rect 784 1283 795 1317
rect 739 1249 795 1283
rect 739 1215 750 1249
rect 784 1215 795 1249
rect 739 1181 795 1215
rect 739 1147 750 1181
rect 784 1147 795 1181
rect 739 1129 795 1147
rect 915 1317 968 1329
rect 915 1283 926 1317
rect 960 1283 968 1317
rect 915 1249 968 1283
rect 915 1215 926 1249
rect 960 1215 968 1249
rect 915 1181 968 1215
rect 915 1147 926 1181
rect 960 1147 968 1181
rect 915 1129 968 1147
rect 1226 930 1279 948
rect 1226 896 1234 930
rect 1268 896 1279 930
rect 1226 862 1279 896
rect 1226 828 1234 862
rect 1268 828 1279 862
rect 1226 794 1279 828
rect 1226 760 1234 794
rect 1268 760 1279 794
rect 1226 748 1279 760
rect 1399 930 1452 948
rect 1399 896 1410 930
rect 1444 896 1452 930
rect 1399 862 1452 896
rect 1399 828 1410 862
rect 1444 828 1452 862
rect 1399 794 1452 828
rect 1399 760 1410 794
rect 1444 760 1452 794
rect 1399 748 1452 760
rect 1226 668 1279 680
rect 1226 634 1234 668
rect 1268 634 1279 668
rect 1226 600 1279 634
rect 1226 566 1234 600
rect 1268 566 1279 600
rect 1226 532 1279 566
rect 1226 498 1234 532
rect 1268 498 1279 532
rect 1226 480 1279 498
rect 1399 668 1452 680
rect 1399 634 1410 668
rect 1444 634 1452 668
rect 1399 600 1452 634
rect 1399 566 1410 600
rect 1444 566 1452 600
rect 1399 532 1452 566
rect 1399 498 1410 532
rect 1444 498 1452 532
rect 1399 480 1452 498
rect 24771 -1311 24824 -1293
rect 24771 -1345 24779 -1311
rect 24813 -1345 24824 -1311
rect 24771 -1379 24824 -1345
rect 24771 -1413 24779 -1379
rect 24813 -1413 24824 -1379
rect 24771 -1447 24824 -1413
rect 24771 -1481 24779 -1447
rect 24813 -1481 24824 -1447
rect 24771 -1493 24824 -1481
rect 24944 -1379 25000 -1293
rect 24944 -1413 24955 -1379
rect 24989 -1413 25000 -1379
rect 24944 -1447 25000 -1413
rect 24944 -1481 24955 -1447
rect 24989 -1481 25000 -1447
rect 24944 -1493 25000 -1481
rect 25120 -1311 25173 -1293
rect 25120 -1345 25131 -1311
rect 25165 -1345 25173 -1311
rect 25120 -1379 25173 -1345
rect 25120 -1413 25131 -1379
rect 25165 -1413 25173 -1379
rect 25120 -1447 25173 -1413
rect 25120 -1481 25131 -1447
rect 25165 -1481 25173 -1447
rect 25120 -1493 25173 -1481
rect 24771 -1573 24824 -1561
rect 24771 -1607 24779 -1573
rect 24813 -1607 24824 -1573
rect 24771 -1641 24824 -1607
rect 24771 -1675 24779 -1641
rect 24813 -1675 24824 -1641
rect 24771 -1709 24824 -1675
rect 24771 -1743 24779 -1709
rect 24813 -1743 24824 -1709
rect 24771 -1761 24824 -1743
rect 24944 -1573 25000 -1561
rect 24944 -1607 24955 -1573
rect 24989 -1607 25000 -1573
rect 24944 -1641 25000 -1607
rect 24944 -1675 24955 -1641
rect 24989 -1675 25000 -1641
rect 24944 -1709 25000 -1675
rect 24944 -1743 24955 -1709
rect 24989 -1743 25000 -1709
rect 24944 -1761 25000 -1743
rect 25120 -1573 25173 -1561
rect 25120 -1607 25131 -1573
rect 25165 -1607 25173 -1573
rect 25120 -1641 25173 -1607
rect 25120 -1675 25131 -1641
rect 25165 -1675 25173 -1641
rect 25120 -1709 25173 -1675
rect 25120 -1743 25131 -1709
rect 25165 -1743 25173 -1709
rect 25120 -1761 25173 -1743
<< ndiffc >>
rect 1234 236 1268 270
rect 1234 168 1268 202
<< mvndiffc >>
rect 288 1875 322 1909
rect 288 1807 322 1841
rect 464 1875 498 1909
rect 464 1807 498 1841
rect 574 1875 608 1909
rect 574 1807 608 1841
rect 926 1875 960 1909
rect 926 1807 960 1841
rect 1410 236 1444 270
rect 1410 168 1444 202
rect 24779 -1015 24813 -981
rect 24779 -1083 24813 -1049
rect 24955 -1015 24989 -981
rect 24955 -1083 24989 -1049
rect 25131 -1015 25165 -981
rect 25131 -1083 25165 -1049
<< mvpdiffc >>
rect 288 1545 322 1579
rect 288 1477 322 1511
rect 288 1409 322 1443
rect 464 1545 498 1579
rect 464 1477 498 1511
rect 464 1409 498 1443
rect 574 1545 608 1579
rect 574 1477 608 1511
rect 574 1409 608 1443
rect 750 1545 784 1579
rect 750 1477 784 1511
rect 750 1409 784 1443
rect 926 1545 960 1579
rect 926 1477 960 1511
rect 926 1409 960 1443
rect 288 1283 322 1317
rect 288 1215 322 1249
rect 288 1147 322 1181
rect 464 1283 498 1317
rect 464 1215 498 1249
rect 464 1147 498 1181
rect 574 1283 608 1317
rect 574 1215 608 1249
rect 574 1147 608 1181
rect 750 1283 784 1317
rect 750 1215 784 1249
rect 750 1147 784 1181
rect 926 1283 960 1317
rect 926 1215 960 1249
rect 926 1147 960 1181
rect 1234 896 1268 930
rect 1234 828 1268 862
rect 1234 760 1268 794
rect 1410 896 1444 930
rect 1410 828 1444 862
rect 1410 760 1444 794
rect 1234 634 1268 668
rect 1234 566 1268 600
rect 1234 498 1268 532
rect 1410 634 1444 668
rect 1410 566 1444 600
rect 1410 498 1444 532
rect 24779 -1345 24813 -1311
rect 24779 -1413 24813 -1379
rect 24779 -1481 24813 -1447
rect 24955 -1413 24989 -1379
rect 24955 -1481 24989 -1447
rect 25131 -1345 25165 -1311
rect 25131 -1413 25165 -1379
rect 25131 -1481 25165 -1447
rect 24779 -1607 24813 -1573
rect 24779 -1675 24813 -1641
rect 24779 -1743 24813 -1709
rect 24955 -1607 24989 -1573
rect 24955 -1675 24989 -1641
rect 24955 -1743 24989 -1709
rect 25131 -1607 25165 -1573
rect 25131 -1675 25165 -1641
rect 25131 -1743 25165 -1709
<< mvpsubdiff >>
rect 265 2010 299 2044
rect 333 2010 390 2044
rect 424 2010 481 2044
rect 515 2010 572 2044
rect 606 2010 663 2044
rect 697 2010 754 2044
rect 788 2010 845 2044
rect 879 2010 939 2044
rect 281 33 315 67
rect 349 33 457 67
rect 491 33 600 67
rect 634 33 743 67
rect 777 33 886 67
rect 920 33 1029 67
rect 1063 33 1172 67
rect 1206 33 1315 67
rect 1349 33 1458 67
rect 1492 33 1526 67
<< mvnsubdiff >>
rect 245 1022 279 1056
rect 313 1022 349 1056
rect 383 1022 419 1056
rect 453 1022 489 1056
rect 523 1022 559 1056
rect 593 1022 629 1056
rect 663 1022 699 1056
rect 733 1022 769 1056
rect 803 1022 839 1056
rect 873 1022 909 1056
rect 943 1022 979 1056
rect 1013 1022 1049 1056
rect 1083 1022 1119 1056
rect 1153 1022 1188 1056
rect 1222 1022 1257 1056
rect 1291 1022 1326 1056
rect 1360 1022 1395 1056
rect 1429 1022 1464 1056
rect 1498 1022 1532 1056
<< mvpsubdiffcont >>
rect 299 2010 333 2044
rect 390 2010 424 2044
rect 481 2010 515 2044
rect 572 2010 606 2044
rect 663 2010 697 2044
rect 754 2010 788 2044
rect 845 2010 879 2044
rect 315 33 349 67
rect 457 33 491 67
rect 600 33 634 67
rect 743 33 777 67
rect 886 33 920 67
rect 1029 33 1063 67
rect 1172 33 1206 67
rect 1315 33 1349 67
rect 1458 33 1492 67
<< mvnsubdiffcont >>
rect 279 1022 313 1056
rect 349 1022 383 1056
rect 419 1022 453 1056
rect 489 1022 523 1056
rect 559 1022 593 1056
rect 629 1022 663 1056
rect 699 1022 733 1056
rect 769 1022 803 1056
rect 839 1022 873 1056
rect 909 1022 943 1056
rect 979 1022 1013 1056
rect 1049 1022 1083 1056
rect 1119 1022 1153 1056
rect 1188 1022 1222 1056
rect 1257 1022 1291 1056
rect 1326 1022 1360 1056
rect 1395 1022 1429 1056
rect 1464 1022 1498 1056
<< poly >>
rect 333 1935 453 1961
rect 619 1935 739 1961
rect 795 1935 915 1961
rect 333 1747 453 1795
rect 333 1713 375 1747
rect 409 1713 453 1747
rect 333 1679 453 1713
rect 333 1645 375 1679
rect 409 1645 453 1679
rect 333 1597 453 1645
rect 619 1747 739 1795
rect 619 1713 664 1747
rect 698 1713 739 1747
rect 619 1679 739 1713
rect 619 1645 664 1679
rect 698 1645 739 1679
rect 619 1597 739 1645
rect 795 1747 915 1795
rect 795 1713 835 1747
rect 869 1713 915 1747
rect 795 1679 915 1713
rect 795 1645 835 1679
rect 869 1645 915 1679
rect 795 1597 915 1645
rect 333 1329 453 1397
rect 619 1329 739 1397
rect 795 1329 915 1397
rect 333 1103 453 1129
rect 619 1103 739 1129
rect 795 1103 915 1129
rect 1279 948 1399 974
rect 1279 680 1399 748
rect 1279 432 1399 480
rect 1279 398 1323 432
rect 1357 398 1399 432
rect 1279 364 1399 398
rect 1279 330 1323 364
rect 1357 330 1399 364
rect 1279 282 1399 330
rect 1279 116 1399 142
rect 24824 -955 24944 -929
rect 25000 -955 25120 -929
rect 24824 -1143 24944 -1095
rect 24824 -1177 24867 -1143
rect 24901 -1177 24944 -1143
rect 24824 -1211 24944 -1177
rect 24824 -1245 24867 -1211
rect 24901 -1245 24944 -1211
rect 24824 -1293 24944 -1245
rect 25000 -1143 25120 -1095
rect 25000 -1177 25045 -1143
rect 25079 -1177 25120 -1143
rect 25000 -1211 25120 -1177
rect 25000 -1245 25045 -1211
rect 25079 -1245 25120 -1211
rect 25000 -1293 25120 -1245
rect 24824 -1561 24944 -1493
rect 25000 -1561 25120 -1493
rect 24824 -1787 24944 -1761
rect 25000 -1787 25120 -1761
<< polycont >>
rect 375 1713 409 1747
rect 375 1645 409 1679
rect 664 1713 698 1747
rect 664 1645 698 1679
rect 835 1713 869 1747
rect 835 1645 869 1679
rect 1323 398 1357 432
rect 1323 330 1357 364
rect 24867 -1177 24901 -1143
rect 24867 -1245 24901 -1211
rect 25045 -1177 25079 -1143
rect 25045 -1245 25079 -1211
<< locali >>
rect 285 2044 323 2049
rect 357 2044 395 2049
rect 285 2015 299 2044
rect 357 2015 390 2044
rect 429 2015 467 2049
rect 501 2044 539 2049
rect 573 2044 611 2049
rect 515 2015 539 2044
rect 606 2015 611 2044
rect 645 2044 683 2049
rect 717 2044 755 2049
rect 645 2015 663 2044
rect 717 2015 754 2044
rect 789 2015 827 2049
rect 265 2010 299 2015
rect 333 2010 390 2015
rect 424 2010 481 2015
rect 515 2010 572 2015
rect 606 2010 663 2015
rect 697 2010 754 2015
rect 788 2010 845 2015
rect 879 2010 913 2044
rect 288 1909 322 1925
rect 288 1841 322 1875
rect 288 1680 322 1807
rect 464 1909 498 1924
rect 464 1841 498 1852
rect 464 1791 498 1807
rect 574 1909 613 1925
rect 608 1875 613 1909
rect 574 1852 613 1875
rect 926 1909 960 1924
rect 574 1841 784 1852
rect 608 1818 784 1841
rect 574 1791 608 1807
rect 288 1608 322 1646
rect 359 1713 375 1747
rect 409 1713 431 1714
rect 359 1679 431 1713
rect 359 1645 375 1679
rect 409 1676 431 1679
rect 648 1713 664 1747
rect 698 1713 714 1714
rect 648 1679 714 1713
rect 648 1645 664 1679
rect 698 1676 714 1679
rect 288 1511 322 1545
rect 288 1443 322 1477
rect 288 1317 322 1409
rect 288 1249 322 1283
rect 288 1181 322 1215
rect 288 1129 322 1147
rect 464 1579 498 1595
rect 464 1511 498 1545
rect 464 1443 498 1477
rect 464 1317 498 1409
rect 464 1249 498 1283
rect 464 1207 498 1215
rect 464 1135 498 1147
rect 574 1579 608 1595
rect 574 1511 608 1545
rect 574 1443 608 1477
rect 574 1317 608 1409
rect 574 1249 608 1283
rect 574 1207 608 1215
rect 574 1135 608 1147
rect 750 1579 784 1818
rect 926 1841 960 1852
rect 926 1791 960 1807
rect 819 1713 835 1747
rect 869 1713 891 1714
rect 819 1679 891 1713
rect 819 1645 835 1679
rect 869 1676 891 1679
rect 750 1511 784 1545
rect 926 1579 960 1595
rect 926 1511 960 1545
rect 750 1476 756 1477
rect 750 1443 790 1476
rect 784 1438 790 1443
rect 750 1404 756 1409
rect 926 1443 960 1477
rect 750 1317 784 1404
rect 750 1249 784 1283
rect 750 1181 784 1215
rect 750 1129 784 1147
rect 926 1317 960 1409
rect 926 1249 960 1283
rect 926 1207 960 1215
rect 926 1135 960 1147
rect 219 1028 259 1062
rect 293 1056 333 1062
rect 367 1056 407 1062
rect 441 1056 481 1062
rect 515 1056 555 1062
rect 589 1056 629 1062
rect 663 1056 703 1062
rect 737 1056 777 1062
rect 811 1056 851 1062
rect 885 1056 925 1062
rect 959 1056 999 1062
rect 1033 1056 1073 1062
rect 1107 1056 1147 1062
rect 1181 1056 1221 1062
rect 1255 1056 1296 1062
rect 1330 1056 1371 1062
rect 1405 1056 1446 1062
rect 1480 1056 1521 1062
rect 313 1028 333 1056
rect 383 1028 407 1056
rect 453 1028 481 1056
rect 523 1028 555 1056
rect 245 1022 279 1028
rect 313 1022 349 1028
rect 383 1022 419 1028
rect 453 1022 489 1028
rect 523 1022 559 1028
rect 593 1022 629 1056
rect 663 1022 699 1056
rect 737 1028 769 1056
rect 811 1028 839 1056
rect 885 1028 909 1056
rect 959 1028 979 1056
rect 1033 1028 1049 1056
rect 1107 1028 1119 1056
rect 1181 1028 1188 1056
rect 1255 1028 1257 1056
rect 733 1022 769 1028
rect 803 1022 839 1028
rect 873 1022 909 1028
rect 943 1022 979 1028
rect 1013 1022 1049 1028
rect 1083 1022 1119 1028
rect 1153 1022 1188 1028
rect 1222 1022 1257 1028
rect 1291 1028 1296 1056
rect 1360 1028 1371 1056
rect 1429 1028 1446 1056
rect 1498 1028 1521 1056
rect 1555 1028 1596 1062
rect 1291 1022 1326 1028
rect 1360 1022 1395 1028
rect 1429 1022 1464 1028
rect 1498 1022 1532 1028
rect 1234 930 1268 942
rect 1234 862 1268 870
rect 1234 794 1268 828
rect 1234 668 1268 760
rect 1234 600 1268 634
rect 1410 930 1444 948
rect 1410 862 1444 896
rect 1410 794 1444 828
rect 1410 668 1444 760
rect 1410 632 1444 634
rect 1360 598 1398 632
rect 1432 600 1444 632
rect 1234 532 1268 566
rect 1234 482 1268 498
rect 1410 532 1444 566
rect 1307 401 1319 432
rect 1307 398 1323 401
rect 1357 398 1373 432
rect 1307 364 1373 398
rect 1307 363 1323 364
rect 1307 330 1319 363
rect 1357 330 1373 364
rect 1234 225 1268 286
rect 1234 153 1268 191
rect 1410 270 1444 498
rect 1410 202 1444 236
rect 1410 152 1444 168
rect 281 33 315 67
rect 349 33 457 67
rect 491 66 600 67
rect 634 66 743 67
rect 777 66 886 67
rect 920 66 1029 67
rect 1063 66 1172 67
rect 1206 66 1315 67
rect 1349 66 1458 67
rect 491 33 568 66
rect 634 33 642 66
rect 602 32 642 33
rect 676 32 716 66
rect 777 33 789 66
rect 750 32 789 33
rect 823 32 862 66
rect 920 33 935 66
rect 896 32 935 33
rect 969 32 1008 66
rect 1063 33 1081 66
rect 1042 32 1081 33
rect 1115 32 1154 66
rect 1206 33 1227 66
rect 1188 32 1227 33
rect 1261 32 1300 66
rect 1349 33 1373 66
rect 1334 32 1373 33
rect 1407 32 1446 66
rect 1492 33 1526 67
rect 24779 -981 24813 -966
rect 24779 -1049 24813 -1038
rect 24779 -1099 24813 -1083
rect 24955 -981 24989 -965
rect 24955 -1049 24989 -1015
rect 24851 -1189 24867 -1143
rect 24901 -1189 24917 -1143
rect 24851 -1211 24917 -1189
rect 24851 -1245 24867 -1211
rect 24901 -1245 24917 -1211
rect 24955 -1295 24989 -1083
rect 25131 -981 25165 -966
rect 25131 -1049 25165 -1038
rect 25131 -1099 25165 -1083
rect 25029 -1189 25045 -1143
rect 25079 -1189 25095 -1143
rect 25029 -1211 25095 -1189
rect 25029 -1245 25045 -1211
rect 25079 -1245 25095 -1211
rect 24779 -1311 24813 -1295
rect 24955 -1307 25165 -1295
rect 24955 -1329 25131 -1307
rect 24779 -1379 24813 -1345
rect 24779 -1447 24813 -1413
rect 24779 -1573 24813 -1481
rect 24779 -1641 24813 -1607
rect 24779 -1683 24813 -1675
rect 24779 -1755 24813 -1743
rect 24955 -1379 24989 -1363
rect 24955 -1447 24989 -1413
rect 24955 -1573 24989 -1481
rect 24955 -1641 24989 -1607
rect 24955 -1709 24989 -1675
rect 24955 -1759 24989 -1743
rect 25131 -1379 25165 -1345
rect 25131 -1447 25165 -1413
rect 25131 -1573 25165 -1481
rect 25131 -1641 25165 -1607
rect 25131 -1709 25165 -1675
rect 25131 -1789 25165 -1743
<< viali >>
rect 251 2015 285 2049
rect 323 2044 357 2049
rect 395 2044 429 2049
rect 323 2015 333 2044
rect 333 2015 357 2044
rect 395 2015 424 2044
rect 424 2015 429 2044
rect 467 2044 501 2049
rect 539 2044 573 2049
rect 467 2015 481 2044
rect 481 2015 501 2044
rect 539 2015 572 2044
rect 572 2015 573 2044
rect 611 2015 645 2049
rect 683 2044 717 2049
rect 755 2044 789 2049
rect 683 2015 697 2044
rect 697 2015 717 2044
rect 755 2015 788 2044
rect 788 2015 789 2044
rect 827 2044 861 2049
rect 827 2015 845 2044
rect 845 2015 861 2044
rect 464 1924 498 1958
rect 464 1875 498 1886
rect 464 1852 498 1875
rect 926 1924 960 1958
rect 926 1875 960 1886
rect 926 1852 960 1875
rect 397 1747 431 1748
rect 680 1747 714 1748
rect 288 1646 322 1680
rect 397 1714 409 1747
rect 409 1714 431 1747
rect 397 1645 409 1676
rect 409 1645 431 1676
rect 680 1714 698 1747
rect 698 1714 714 1747
rect 680 1645 698 1676
rect 698 1645 714 1676
rect 397 1642 431 1645
rect 680 1642 714 1645
rect 288 1579 322 1608
rect 288 1574 322 1579
rect 464 1181 498 1207
rect 464 1173 498 1181
rect 464 1101 498 1135
rect 574 1181 608 1207
rect 574 1173 608 1181
rect 574 1101 608 1135
rect 857 1747 891 1748
rect 857 1714 869 1747
rect 869 1714 891 1747
rect 857 1645 869 1676
rect 869 1645 891 1676
rect 857 1642 891 1645
rect 756 1477 784 1510
rect 784 1477 790 1510
rect 756 1476 790 1477
rect 756 1409 784 1438
rect 784 1409 790 1438
rect 756 1404 790 1409
rect 926 1181 960 1207
rect 926 1173 960 1181
rect 926 1101 960 1135
rect 185 1028 219 1062
rect 259 1056 293 1062
rect 333 1056 367 1062
rect 407 1056 441 1062
rect 481 1056 515 1062
rect 555 1056 589 1062
rect 629 1056 663 1062
rect 703 1056 737 1062
rect 777 1056 811 1062
rect 851 1056 885 1062
rect 925 1056 959 1062
rect 999 1056 1033 1062
rect 1073 1056 1107 1062
rect 1147 1056 1181 1062
rect 1221 1056 1255 1062
rect 1296 1056 1330 1062
rect 1371 1056 1405 1062
rect 1446 1056 1480 1062
rect 259 1028 279 1056
rect 279 1028 293 1056
rect 333 1028 349 1056
rect 349 1028 367 1056
rect 407 1028 419 1056
rect 419 1028 441 1056
rect 481 1028 489 1056
rect 489 1028 515 1056
rect 555 1028 559 1056
rect 559 1028 589 1056
rect 629 1028 663 1056
rect 703 1028 733 1056
rect 733 1028 737 1056
rect 777 1028 803 1056
rect 803 1028 811 1056
rect 851 1028 873 1056
rect 873 1028 885 1056
rect 925 1028 943 1056
rect 943 1028 959 1056
rect 999 1028 1013 1056
rect 1013 1028 1033 1056
rect 1073 1028 1083 1056
rect 1083 1028 1107 1056
rect 1147 1028 1153 1056
rect 1153 1028 1181 1056
rect 1221 1028 1222 1056
rect 1222 1028 1255 1056
rect 1296 1028 1326 1056
rect 1326 1028 1330 1056
rect 1371 1028 1395 1056
rect 1395 1028 1405 1056
rect 1446 1028 1464 1056
rect 1464 1028 1480 1056
rect 1521 1028 1555 1062
rect 1596 1028 1630 1062
rect 1234 942 1268 976
rect 1234 896 1268 904
rect 1234 870 1268 896
rect 1326 598 1360 632
rect 1398 600 1432 632
rect 1398 598 1410 600
rect 1410 598 1432 600
rect 1319 432 1353 435
rect 1319 401 1323 432
rect 1323 401 1353 432
rect 1319 330 1323 363
rect 1323 330 1353 363
rect 1319 329 1353 330
rect 1234 191 1268 225
rect 1234 119 1268 153
rect 568 33 600 66
rect 600 33 602 66
rect 568 32 602 33
rect 642 32 676 66
rect 716 33 743 66
rect 743 33 750 66
rect 716 32 750 33
rect 789 32 823 66
rect 862 33 886 66
rect 886 33 896 66
rect 862 32 896 33
rect 935 32 969 66
rect 1008 33 1029 66
rect 1029 33 1042 66
rect 1008 32 1042 33
rect 1081 32 1115 66
rect 1154 33 1172 66
rect 1172 33 1188 66
rect 1154 32 1188 33
rect 1227 32 1261 66
rect 1300 33 1315 66
rect 1315 33 1334 66
rect 1300 32 1334 33
rect 1373 32 1407 66
rect 1446 33 1458 66
rect 1458 33 1480 66
rect 1446 32 1480 33
rect 24779 -966 24813 -932
rect 24779 -1015 24813 -1004
rect 24779 -1038 24813 -1015
rect 24867 -1177 24901 -1155
rect 24867 -1189 24901 -1177
rect 24867 -1245 24901 -1227
rect 24867 -1261 24901 -1245
rect 25131 -966 25165 -932
rect 25131 -1015 25165 -1004
rect 25131 -1038 25165 -1015
rect 25045 -1177 25079 -1155
rect 25045 -1189 25079 -1177
rect 25045 -1245 25079 -1227
rect 25045 -1261 25079 -1245
rect 25131 -1311 25165 -1307
rect 25131 -1341 25165 -1311
rect 24779 -1709 24813 -1683
rect 24779 -1717 24813 -1709
rect 24779 -1789 24813 -1755
rect 25131 -1413 25165 -1379
<< metal1 >>
rect 20418 2665 20424 2717
rect 20476 2665 20488 2717
rect 20540 2665 22488 2717
rect 22540 2665 22552 2717
rect 22604 2665 22610 2717
rect 233 2049 1010 2055
rect 233 2015 251 2049
rect 285 2015 323 2049
rect 357 2015 395 2049
rect 429 2015 467 2049
rect 501 2015 539 2049
rect 573 2015 611 2049
rect 645 2015 683 2049
rect 717 2015 755 2049
rect 789 2015 827 2049
rect 861 2015 1010 2049
rect 233 1958 1010 2015
rect 233 1924 464 1958
rect 498 1924 926 1958
rect 960 1924 1010 1958
rect 233 1886 1010 1924
rect 11109 1913 11446 2058
rect 233 1852 464 1886
rect 498 1852 926 1886
rect 960 1852 1010 1886
rect 233 1840 1010 1852
rect 391 1748 437 1760
rect 391 1714 397 1748
rect 431 1714 437 1748
rect 282 1684 337 1692
rect 282 1632 285 1684
rect 282 1620 337 1632
rect 282 1568 285 1620
rect 282 1562 337 1568
rect 391 1676 437 1714
rect 391 1642 397 1676
rect 431 1642 437 1676
rect 391 1522 437 1642
rect 674 1752 729 1760
rect 674 1700 677 1752
rect 674 1688 729 1700
rect 674 1636 677 1688
rect 674 1630 729 1636
rect 848 1752 900 1760
rect 2391 1754 2470 1760
rect 848 1688 900 1700
rect 2357 1658 2379 1721
rect 2391 1702 2418 1754
rect 2391 1690 2470 1702
rect 848 1630 900 1636
rect 2391 1638 2418 1690
rect 2391 1630 2470 1638
rect 2058 1578 2183 1584
tri 437 1522 471 1556 sw
rect 2110 1526 2183 1578
rect 391 1510 796 1522
rect 391 1476 756 1510
rect 790 1476 796 1510
rect 391 1470 796 1476
tri 716 1438 748 1470 ne
rect 748 1438 796 1470
rect 2058 1514 2183 1526
rect 2110 1462 2183 1514
rect 2321 1490 2442 1561
rect 2058 1454 2183 1462
tri 748 1436 750 1438 ne
rect 750 1404 756 1438
rect 790 1404 796 1438
rect 3897 1427 3939 1510
rect 750 1392 796 1404
rect 173 1220 269 1221
rect 173 1207 1009 1220
rect 11163 1208 11555 1356
rect 173 1173 464 1207
rect 498 1173 574 1207
rect 608 1173 926 1207
rect 960 1173 1009 1207
rect 173 1135 1009 1173
rect 173 1101 464 1135
rect 498 1101 574 1135
rect 608 1101 926 1135
rect 960 1101 1009 1135
rect 173 1068 1009 1101
rect 173 1062 1642 1068
rect 173 1028 185 1062
rect 219 1028 259 1062
rect 293 1028 333 1062
rect 367 1028 407 1062
rect 441 1028 481 1062
rect 515 1028 555 1062
rect 589 1028 629 1062
rect 663 1028 703 1062
rect 737 1028 777 1062
rect 811 1028 851 1062
rect 885 1028 925 1062
rect 959 1028 999 1062
rect 1033 1028 1073 1062
rect 1107 1028 1147 1062
rect 1181 1028 1221 1062
rect 1255 1028 1296 1062
rect 1330 1028 1371 1062
rect 1405 1028 1446 1062
rect 1480 1028 1521 1062
rect 1555 1028 1596 1062
rect 1630 1060 1642 1062
rect 1630 1028 1672 1060
rect 173 1022 1672 1028
rect 173 1017 1009 1022
rect 173 857 879 1017
rect 1104 976 1672 1022
rect 1104 942 1234 976
rect 1268 942 1672 976
rect 1104 904 1672 942
rect 1104 870 1234 904
rect 1268 870 1672 904
rect 1104 858 1672 870
rect 1179 857 1499 858
rect 4979 735 4985 787
rect 5037 735 5049 787
rect 5101 735 5107 787
rect 1201 716 1253 722
rect 1067 704 1119 705
rect 974 699 1119 704
rect 974 658 1067 699
rect 1067 635 1119 647
rect 1201 650 1253 664
rect 1924 643 1988 695
rect 2040 643 2052 695
rect 2104 643 2629 695
rect 2681 643 2693 695
rect 2745 643 2751 695
rect 1253 632 1444 638
rect 1253 598 1326 632
rect 1360 598 1398 632
rect 1432 598 1444 632
rect 1201 592 1444 598
rect 1067 577 1119 583
rect 1313 435 1359 447
rect 1313 401 1319 435
rect 1353 401 1359 435
rect 1143 357 1282 393
rect 1313 363 1359 401
rect 1313 329 1319 363
rect 1353 329 1359 363
rect 1313 317 1359 329
rect 3413 397 3465 403
rect 3413 333 3465 345
rect 3413 275 3465 281
rect 804 72 879 237
rect 1180 225 1574 237
rect 1180 191 1234 225
rect 1268 191 1574 225
rect 10997 211 11468 379
rect 1180 153 1574 191
rect 1180 119 1234 153
rect 1268 119 1574 153
rect 1180 72 1574 119
rect 556 66 1574 72
rect 556 32 568 66
rect 602 32 642 66
rect 676 32 716 66
rect 750 32 789 66
rect 823 32 862 66
rect 896 32 935 66
rect 969 32 1008 66
rect 1042 32 1081 66
rect 1115 32 1154 66
rect 1188 32 1227 66
rect 1261 32 1300 66
rect 1334 32 1373 66
rect 1407 32 1446 66
rect 1480 32 1574 66
rect 556 26 1574 32
rect 804 23 879 26
rect 1180 23 1574 26
rect 1180 22 1499 23
tri 4517 -11 4525 -3 se
rect 4525 -11 16541 -3
rect 1319 -63 3378 -11
rect 3430 -63 3442 -11
rect 3494 -55 16541 -11
rect 3494 -63 4539 -55
tri 4539 -63 4547 -55 nw
rect 12604 -135 20056 -83
rect 20108 -135 20120 -83
rect 20172 -135 20178 -83
tri 2633 -407 2685 -355 se
rect 2685 -407 22131 -355
rect 22183 -407 22195 -355
rect 22247 -407 22253 -355
tri 2611 -429 2633 -407 se
rect 2633 -429 2685 -407
tri 2685 -429 2707 -407 nw
tri 2537 -503 2611 -429 se
tri 2611 -503 2685 -429 nw
rect 20655 -487 20661 -435
rect 20713 -487 20725 -435
rect 20777 -487 22262 -435
rect 22314 -487 22326 -435
rect 22378 -487 22384 -435
tri 2463 -577 2537 -503 se
tri 2537 -577 2611 -503 nw
rect 22900 -567 22906 -515
rect 22958 -567 22970 -515
rect 23022 -567 24859 -515
rect 24911 -567 24923 -515
rect 24975 -567 24990 -515
tri 2389 -651 2463 -577 se
tri 2463 -651 2537 -577 nw
tri 2335 -705 2389 -651 se
rect 2389 -705 2409 -651
tri 2409 -705 2463 -651 nw
rect 543 -757 553 -705
rect 605 -757 617 -705
rect 669 -757 2357 -705
tri 2357 -757 2409 -705 nw
rect 22340 -807 22346 -755
rect 22398 -807 22410 -755
rect 22462 -807 24688 -755
rect 24740 -807 24752 -755
rect 24804 -807 24810 -755
rect 24746 -932 25177 -835
rect 24746 -966 24779 -932
rect 24813 -966 25131 -932
rect 25165 -966 25177 -932
rect 24746 -1004 25177 -966
rect 24746 -1038 24779 -1004
rect 24813 -1038 25131 -1004
rect 25165 -1038 25177 -1004
rect 24746 -1050 25177 -1038
rect 24851 -1149 24907 -1143
rect 24903 -1201 24907 -1149
rect 24851 -1215 24907 -1201
rect 24903 -1267 24907 -1215
rect 24851 -1273 24907 -1267
rect 25036 -1149 25088 -1143
rect 25036 -1215 25088 -1201
rect 25036 -1273 25088 -1267
rect 25122 -1301 25174 -1295
rect 25122 -1367 25174 -1353
rect 25122 -1425 25174 -1419
rect 24767 -1683 25177 -1670
rect 24767 -1717 24779 -1683
rect 24813 -1717 25177 -1683
rect 24767 -1755 25177 -1717
rect 24767 -1789 24779 -1755
rect 24813 -1789 25177 -1755
rect 24767 -1873 25177 -1789
<< via1 >>
rect 20424 2665 20476 2717
rect 20488 2665 20540 2717
rect 22488 2665 22540 2717
rect 22552 2665 22604 2717
rect 285 1680 337 1684
rect 285 1646 288 1680
rect 288 1646 322 1680
rect 322 1646 337 1680
rect 285 1632 337 1646
rect 285 1608 337 1620
rect 285 1574 288 1608
rect 288 1574 322 1608
rect 322 1574 337 1608
rect 285 1568 337 1574
rect 677 1748 729 1752
rect 677 1714 680 1748
rect 680 1714 714 1748
rect 714 1714 729 1748
rect 677 1700 729 1714
rect 677 1676 729 1688
rect 677 1642 680 1676
rect 680 1642 714 1676
rect 714 1642 729 1676
rect 677 1636 729 1642
rect 848 1748 900 1752
rect 848 1714 857 1748
rect 857 1714 891 1748
rect 891 1714 900 1748
rect 848 1700 900 1714
rect 848 1676 900 1688
rect 848 1642 857 1676
rect 857 1642 891 1676
rect 891 1642 900 1676
rect 2418 1702 2470 1754
rect 848 1636 900 1642
rect 2418 1638 2470 1690
rect 2058 1526 2110 1578
rect 2058 1462 2110 1514
rect 4985 735 5037 787
rect 5049 735 5101 787
rect 1067 647 1119 699
rect 1067 583 1119 635
rect 1201 664 1253 716
rect 1201 598 1253 650
rect 1988 643 2040 695
rect 2052 643 2104 695
rect 2629 643 2681 695
rect 2693 643 2745 695
rect 3413 345 3465 397
rect 3413 281 3465 333
rect 3378 -63 3430 -11
rect 3442 -63 3494 -11
rect 20056 -135 20108 -83
rect 20120 -135 20172 -83
rect 22131 -407 22183 -355
rect 22195 -407 22247 -355
rect 20661 -487 20713 -435
rect 20725 -487 20777 -435
rect 22262 -487 22314 -435
rect 22326 -487 22378 -435
rect 22906 -567 22958 -515
rect 22970 -567 23022 -515
rect 24859 -567 24911 -515
rect 24923 -567 24975 -515
rect 553 -757 605 -705
rect 617 -757 669 -705
rect 22346 -807 22398 -755
rect 22410 -807 22462 -755
rect 24688 -807 24740 -755
rect 24752 -807 24804 -755
rect 24851 -1155 24903 -1149
rect 24851 -1189 24867 -1155
rect 24867 -1189 24901 -1155
rect 24901 -1189 24903 -1155
rect 24851 -1201 24903 -1189
rect 24851 -1227 24903 -1215
rect 24851 -1261 24867 -1227
rect 24867 -1261 24901 -1227
rect 24901 -1261 24903 -1227
rect 24851 -1267 24903 -1261
rect 25036 -1155 25088 -1149
rect 25036 -1189 25045 -1155
rect 25045 -1189 25079 -1155
rect 25079 -1189 25088 -1155
rect 25036 -1201 25088 -1189
rect 25036 -1227 25088 -1215
rect 25036 -1261 25045 -1227
rect 25045 -1261 25079 -1227
rect 25079 -1261 25088 -1227
rect 25036 -1267 25088 -1261
rect 25122 -1307 25174 -1301
rect 25122 -1341 25131 -1307
rect 25131 -1341 25165 -1307
rect 25165 -1341 25174 -1307
rect 25122 -1353 25174 -1341
rect 25122 -1379 25174 -1367
rect 25122 -1413 25131 -1379
rect 25131 -1413 25165 -1379
rect 25165 -1413 25174 -1379
rect 25122 -1419 25174 -1413
<< metal2 >>
tri 20363 2665 20415 2717 se
rect 20415 2665 20424 2717
rect 20476 2665 20488 2717
rect 20540 2665 20546 2717
rect 22482 2665 22488 2717
rect 22540 2665 22552 2717
rect 22604 2665 22610 2717
tri 20342 2644 20363 2665 se
rect 20363 2644 20415 2665
tri 20415 2644 20436 2665 nw
tri 20269 2571 20342 2644 se
tri 20342 2571 20415 2644 nw
tri 20251 2553 20269 2571 se
rect 20269 2553 20324 2571
tri 20324 2553 20342 2571 nw
tri 10252 2492 10313 2553 se
rect 10313 2512 20283 2553
tri 20283 2512 20324 2553 nw
tri 10313 2492 10333 2512 nw
tri 10191 2431 10252 2492 se
tri 10252 2431 10313 2492 nw
rect 20131 2431 20305 2443
tri 20305 2431 20317 2443 sw
tri 10130 2370 10191 2431 se
tri 10191 2370 10252 2431 nw
rect 20131 2405 20317 2431
tri 20317 2405 20343 2431 sw
rect 20131 2402 20343 2405
tri 20266 2370 20298 2402 ne
rect 20298 2370 20343 2402
tri 20343 2370 20378 2405 sw
tri 10095 2335 10130 2370 se
rect 10130 2335 10156 2370
tri 10156 2335 10191 2370 nw
tri 20298 2335 20333 2370 ne
rect 20333 2335 20378 2370
tri 20378 2335 20413 2370 sw
rect 3995 2294 4013 2335
rect 4004 2279 4013 2294
rect 4069 2279 4093 2335
rect 4149 2294 10115 2335
tri 10115 2294 10156 2335 nw
tri 20333 2325 20343 2335 ne
rect 20343 2325 20413 2335
tri 20413 2325 20423 2335 sw
tri 20343 2294 20374 2325 ne
rect 20374 2294 20423 2325
tri 20423 2294 20454 2325 sw
rect 4149 2279 4158 2294
tri 20374 2279 20389 2294 ne
rect 20389 2279 20454 2294
tri 20454 2279 20469 2294 sw
tri 20389 2245 20423 2279 ne
rect 20423 2245 20469 2279
tri 20469 2245 20503 2279 sw
tri 20423 2165 20503 2245 ne
tri 20503 2165 20583 2245 sw
rect 22482 2175 22610 2665
tri 22610 2175 22650 2215 sw
tri 20503 2135 20533 2165 ne
rect 20533 2135 22187 2165
rect 22482 2135 22853 2175
tri 20533 2124 20544 2135 ne
rect 20544 2124 22187 2135
tri 22754 2124 22765 2135 ne
rect 22765 2124 22853 2135
tri 22765 2095 22794 2124 ne
rect 677 1752 729 1758
rect 285 1684 337 1690
rect 285 1620 337 1632
rect 285 661 337 1568
rect 677 1688 729 1700
rect 677 1526 729 1636
rect 848 1752 900 1758
rect 2418 1754 2470 1760
rect 848 1690 900 1700
tri 900 1690 912 1702 sw
rect 2418 1690 2470 1702
rect 848 1688 912 1690
rect 900 1668 912 1688
tri 912 1668 934 1690 sw
rect 900 1644 1007 1668
tri 1007 1644 1031 1668 sw
rect 900 1638 1031 1644
tri 1031 1638 1037 1644 sw
rect 900 1636 1037 1638
rect 848 1616 1037 1636
tri 985 1578 1023 1616 ne
rect 1023 1578 1037 1616
tri 1037 1578 1097 1638 sw
rect 2058 1578 2110 1584
tri 1023 1570 1031 1578 ne
rect 1031 1570 1097 1578
tri 1097 1570 1105 1578 sw
tri 1031 1554 1047 1570 ne
rect 1047 1554 1105 1570
tri 729 1526 757 1554 sw
tri 1047 1526 1075 1554 ne
rect 1075 1526 1105 1554
tri 1105 1526 1149 1570 sw
rect 677 1518 757 1526
tri 757 1518 765 1526 sw
tri 1075 1518 1083 1526 ne
rect 1083 1518 1149 1526
rect 677 1516 948 1518
tri 677 1514 679 1516 ne
rect 679 1514 948 1516
tri 948 1514 952 1518 sw
tri 1083 1514 1087 1518 ne
rect 1087 1514 1149 1518
tri 1149 1514 1161 1526 sw
rect 2058 1514 2110 1526
tri 679 1495 698 1514 ne
rect 698 1496 952 1514
tri 952 1496 970 1514 sw
tri 1087 1496 1105 1514 ne
rect 1105 1496 1161 1514
tri 1161 1496 1179 1514 sw
rect 698 1495 970 1496
tri 970 1495 971 1496 sw
tri 1105 1495 1106 1496 ne
rect 1106 1495 1179 1496
tri 698 1466 727 1495 ne
rect 727 1466 971 1495
tri 926 1462 930 1466 ne
rect 930 1462 971 1466
tri 971 1462 1004 1495 sw
tri 1106 1462 1139 1495 ne
rect 1139 1462 1179 1495
tri 1179 1462 1213 1496 sw
tri 930 1421 971 1462 ne
rect 971 1422 1004 1462
tri 1004 1422 1044 1462 sw
tri 1139 1422 1179 1462 ne
rect 1179 1422 1213 1462
tri 1213 1422 1253 1462 sw
rect 971 1421 1044 1422
tri 1044 1421 1045 1422 sw
tri 1179 1421 1180 1422 ne
rect 1180 1421 1253 1422
tri 971 1347 1045 1421 ne
tri 1045 1400 1066 1421 sw
tri 1180 1400 1201 1421 ne
rect 1045 1347 1066 1400
tri 1066 1347 1119 1400 sw
tri 1045 1325 1067 1347 ne
rect 1067 699 1119 1347
tri 337 661 359 683 sw
tri 285 647 299 661 ne
rect 299 647 359 661
tri 359 647 373 661 sw
tri 299 635 311 647 ne
rect 311 635 373 647
tri 373 635 385 647 sw
rect 1067 635 1119 647
tri 311 591 355 635 ne
rect 355 591 385 635
tri 385 591 429 635 sw
tri 355 587 359 591 ne
rect 359 587 429 591
tri 429 587 433 591 sw
tri 359 583 363 587 ne
rect 363 583 433 587
tri 433 583 437 587 sw
rect 1201 716 1253 1421
rect 2058 695 2110 1462
rect 1201 650 1253 664
rect 1982 643 1988 695
rect 2040 643 2052 695
rect 2104 643 2110 695
rect 1201 591 1253 598
tri 363 513 433 583 ne
rect 433 513 437 583
tri 437 513 507 583 sw
tri 433 463 483 513 ne
rect 483 477 507 513
tri 507 477 543 513 sw
rect 483 463 543 477
tri 543 463 557 477 sw
tri 483 439 507 463 ne
rect 507 439 557 463
tri 557 439 581 463 sw
tri 507 403 543 439 ne
rect 543 425 581 439
tri 581 425 595 439 sw
rect 543 -705 595 425
tri 1051 -135 1067 -119 se
rect 1067 -135 1119 583
rect 2418 519 2470 1638
rect 22794 958 22853 2124
tri 22853 958 22864 969 sw
rect 22794 922 22864 958
tri 22794 852 22864 922 ne
tri 22864 852 22970 958 sw
tri 22864 816 22900 852 ne
rect 4979 735 4985 787
rect 5037 735 5049 787
rect 5101 735 5107 787
tri 5021 701 5055 735 ne
rect 2623 694 2629 695
rect 2615 638 2624 694
rect 2681 643 2693 695
rect 2745 694 2751 695
rect 2680 638 2704 643
rect 2760 638 2769 694
rect 2418 463 2427 519
rect 2483 463 2507 519
rect 2563 463 2572 519
rect 3413 397 3465 403
rect 3413 333 3465 345
rect 3413 -11 3465 281
rect 5055 0 5107 735
rect 7128 79 7170 193
rect 7423 78 7468 196
rect 8662 86 8707 178
rect 8833 92 8868 185
rect 10071 90 10110 227
rect 10366 88 10404 197
rect 11274 82 11312 192
rect 11572 89 11608 219
rect 12817 94 12848 165
rect 12978 86 13016 180
rect 14216 91 14252 218
rect 14512 88 14550 198
rect 15421 84 15459 169
rect 15720 91 15758 187
rect 16956 83 16993 175
rect 17122 80 17161 165
rect 18654 84 18696 176
rect 19865 85 19904 175
rect 21101 81 21141 161
rect 21268 85 21309 177
rect 22513 90 22546 213
rect 22801 102 22844 196
rect 3372 -63 3378 -11
rect 3430 -63 3442 -11
rect 3494 -63 3500 -11
rect 20050 -83 20178 25
rect 20050 -135 20056 -83
rect 20108 -135 20120 -83
rect 20172 -135 20178 -83
tri 1006 -180 1051 -135 se
rect 1051 -146 1119 -135
rect 1051 -180 1085 -146
tri 1085 -180 1119 -146 nw
rect 1006 -189 1062 -180
tri 1062 -203 1085 -180 nw
rect 1006 -269 1062 -245
rect 1006 -334 1062 -325
tri 20401 -311 20452 -260 se
rect 20452 -310 20649 -260
rect 20452 -311 20495 -310
tri 20495 -311 20496 -310 nw
tri 20625 -311 20626 -310 ne
rect 20626 -311 20649 -310
rect 20401 -316 20490 -311
tri 20490 -316 20495 -311 nw
tri 20626 -316 20631 -311 ne
rect 20631 -316 20649 -311
tri 20649 -316 20705 -260 sw
rect 20401 -334 20472 -316
tri 20472 -334 20490 -316 nw
tri 20631 -334 20649 -316 ne
rect 20649 -334 20705 -316
tri 595 -705 646 -654 sw
rect 543 -757 553 -705
rect 605 -757 617 -705
rect 669 -757 675 -705
tri 20336 -1128 20401 -1063 se
rect 20401 -1086 20451 -334
tri 20451 -355 20472 -334 nw
tri 20649 -340 20655 -334 ne
rect 20655 -435 20705 -334
rect 22125 -407 22131 -355
rect 22183 -407 22195 -355
rect 22247 -407 22253 -355
tri 20705 -435 20733 -407 sw
tri 22133 -435 22161 -407 ne
rect 22161 -435 22219 -407
rect 20655 -487 20661 -435
rect 20713 -487 20725 -435
rect 20777 -487 20783 -435
tri 22161 -441 22167 -435 ne
rect 22167 -863 22219 -435
rect 22256 -487 22262 -435
rect 22314 -487 22326 -435
rect 22378 -487 22384 -435
tri 22312 -515 22340 -487 ne
rect 22340 -755 22384 -487
rect 22900 -515 22970 852
rect 23713 91 23747 182
rect 24016 96 24046 224
rect 25248 88 25283 211
rect 25417 92 25454 199
rect 26656 96 26693 214
rect 26950 95 26988 181
rect 25094 -75 25150 -66
rect 25094 -155 25150 -131
rect 25094 -220 25150 -211
rect 24853 -515 24862 -511
rect 24918 -515 24942 -511
rect 22900 -567 22906 -515
rect 22958 -567 22970 -515
rect 23022 -567 23028 -515
rect 24853 -567 24859 -515
rect 24918 -567 24923 -515
rect 24998 -567 25007 -511
tri 22384 -755 22418 -721 sw
rect 24682 -755 24691 -751
rect 24747 -755 24771 -751
rect 22340 -807 22346 -755
rect 22398 -807 22410 -755
rect 22462 -807 22468 -755
rect 24682 -807 24688 -755
rect 24747 -807 24752 -755
rect 24827 -807 24836 -751
rect 22167 -915 25665 -863
rect 20401 -1128 20409 -1086
tri 20409 -1128 20451 -1086 nw
tri 19389 -1139 19400 -1128 se
rect 19400 -1139 20398 -1128
tri 20398 -1139 20409 -1128 nw
tri 19379 -1149 19389 -1139 se
rect 19389 -1149 20388 -1139
tri 20388 -1149 20398 -1139 nw
rect 24834 -1143 24890 -1139
rect 24834 -1148 24903 -1143
rect 24890 -1149 24903 -1148
tri 19327 -1201 19379 -1149 se
rect 19379 -1179 20358 -1149
tri 20358 -1179 20388 -1149 nw
rect 19379 -1201 19405 -1179
tri 19405 -1201 19427 -1179 nw
tri 19322 -1206 19327 -1201 se
rect 19327 -1206 19400 -1201
tri 19400 -1206 19405 -1201 nw
rect 24890 -1204 24903 -1201
tri 19313 -1215 19322 -1206 se
rect 19322 -1215 19391 -1206
tri 19391 -1215 19400 -1206 nw
rect 24834 -1215 24903 -1204
tri 19301 -1227 19313 -1215 se
rect 19313 -1227 19379 -1215
tri 19379 -1227 19391 -1215 nw
tri 19263 -1797 19301 -1759 se
rect 19301 -1771 19351 -1227
tri 19351 -1255 19379 -1227 nw
rect 24834 -1228 24851 -1215
rect 24890 -1273 24903 -1267
rect 24968 -1148 25088 -1139
rect 25024 -1149 25088 -1148
rect 25024 -1201 25036 -1149
rect 25024 -1204 25088 -1201
rect 24968 -1215 25088 -1204
rect 24968 -1228 25036 -1215
rect 24834 -1293 24890 -1284
rect 25024 -1267 25036 -1228
rect 25024 -1273 25088 -1267
rect 24968 -1293 25024 -1284
tri 25024 -1293 25044 -1273 nw
tri 25116 -1301 25122 -1295 se
rect 25122 -1301 25174 -1295
tri 25110 -1307 25116 -1301 se
rect 25116 -1307 25122 -1301
rect 25094 -1316 25122 -1307
rect 25150 -1367 25174 -1353
rect 25094 -1396 25122 -1372
rect 25150 -1425 25174 -1419
tri 25150 -1449 25174 -1425 nw
rect 25094 -1461 25150 -1452
rect 19301 -1797 19325 -1771
tri 19325 -1797 19351 -1771 nw
tri 17738 -1882 17823 -1797 se
rect 17823 -1854 19268 -1797
tri 19268 -1854 19325 -1797 nw
tri 17823 -1882 17851 -1854 nw
tri 17719 -1901 17738 -1882 se
rect 17738 -1901 17804 -1882
tri 17804 -1901 17823 -1882 nw
tri 16006 -1904 16009 -1901 se
rect 16009 -1904 17801 -1901
tri 17801 -1904 17804 -1901 nw
rect 4850 -1913 17754 -1904
rect 4906 -1951 17754 -1913
tri 17754 -1951 17801 -1904 nw
rect 4906 -1954 16051 -1951
tri 16051 -1954 16054 -1951 nw
rect 4850 -1993 4906 -1969
tri 4906 -2006 4958 -1954 nw
rect 4850 -2058 4906 -2049
rect 4850 -3715 4906 -3706
tri 4790 -3808 4850 -3748 se
rect 4850 -3795 4906 -3771
tri 3382 -3856 3430 -3808 se
rect 3430 -3851 4850 -3808
rect 3430 -3856 4906 -3851
rect 1006 -3865 1062 -3856
tri 3355 -3883 3382 -3856 se
rect 3382 -3860 4906 -3856
rect 3382 -3883 3430 -3860
tri 3430 -3883 3453 -3860 nw
tri 3342 -3896 3355 -3883 se
rect 3355 -3896 3417 -3883
tri 3417 -3896 3430 -3883 nw
rect 1062 -3921 3363 -3896
rect 1006 -3945 3363 -3921
rect 1062 -3950 3363 -3945
tri 3363 -3950 3417 -3896 nw
rect 1006 -4010 1062 -4001
<< via2 >>
rect 4013 2279 4069 2335
rect 4093 2279 4149 2335
rect 2624 643 2629 694
rect 2629 643 2680 694
rect 2704 643 2745 694
rect 2745 643 2760 694
rect 2624 638 2680 643
rect 2704 638 2760 643
rect 2427 463 2483 519
rect 2507 463 2563 519
rect 1006 -245 1062 -189
rect 1006 -325 1062 -269
rect 25094 -131 25150 -75
rect 25094 -211 25150 -155
rect 24862 -515 24918 -511
rect 24942 -515 24998 -511
rect 24862 -567 24911 -515
rect 24911 -567 24918 -515
rect 24942 -567 24975 -515
rect 24975 -567 24998 -515
rect 24691 -755 24747 -751
rect 24771 -755 24827 -751
rect 24691 -807 24740 -755
rect 24740 -807 24747 -755
rect 24771 -807 24804 -755
rect 24804 -807 24827 -755
rect 24834 -1149 24890 -1148
rect 24834 -1201 24851 -1149
rect 24851 -1201 24890 -1149
rect 24834 -1204 24890 -1201
rect 24834 -1267 24851 -1228
rect 24851 -1267 24890 -1228
rect 24834 -1284 24890 -1267
rect 24968 -1204 25024 -1148
rect 24968 -1284 25024 -1228
rect 25094 -1353 25122 -1316
rect 25122 -1353 25150 -1316
rect 25094 -1367 25150 -1353
rect 25094 -1372 25122 -1367
rect 25122 -1372 25150 -1367
rect 25094 -1419 25122 -1396
rect 25122 -1419 25150 -1396
rect 25094 -1452 25150 -1419
rect 4850 -1969 4906 -1913
rect 4850 -2049 4906 -1993
rect 4850 -3771 4906 -3715
rect 4850 -3851 4906 -3795
rect 1006 -3921 1062 -3865
rect 1006 -4001 1062 -3945
<< metal3 >>
rect 4008 2335 4154 2340
rect 4008 2279 4013 2335
rect 4069 2279 4093 2335
rect 4149 2279 4154 2335
rect 4008 2274 4154 2279
rect 4006 699 4072 2274
rect 2613 694 4072 699
rect 2613 638 2624 694
rect 2680 638 2704 694
rect 2760 638 4072 694
rect 2613 633 4072 638
rect 2422 519 3635 524
rect 2422 463 2427 519
rect 2483 463 2507 519
rect 2563 463 3635 519
rect 2422 458 3635 463
rect 1001 -189 1067 -168
rect 1001 -245 1006 -189
rect 1062 -245 1067 -189
rect 1001 -269 1067 -245
rect 1001 -325 1006 -269
rect 1062 -325 1067 -269
rect 1001 -3865 1067 -325
rect 1001 -3921 1006 -3865
rect 1062 -3921 1067 -3865
rect 1001 -3945 1067 -3921
rect 1001 -4001 1006 -3945
rect 1062 -4001 1067 -3945
rect 1001 -4115 1067 -4001
rect 4006 -4115 4072 633
rect 25089 -75 25155 -70
rect 25089 -131 25094 -75
rect 25150 -131 25155 -75
rect 25089 -155 25155 -131
rect 25089 -211 25094 -155
rect 25150 -211 25155 -155
rect 24857 -511 25029 -506
rect 24857 -567 24862 -511
rect 24918 -567 24942 -511
rect 24998 -567 25029 -511
rect 24857 -572 25029 -567
tri 24897 -638 24963 -572 ne
rect 24673 -751 24868 -746
rect 24673 -807 24691 -751
rect 24747 -807 24771 -751
rect 24827 -773 24868 -751
tri 24868 -773 24895 -746 sw
rect 24827 -807 24895 -773
rect 24673 -812 24895 -807
tri 24799 -842 24829 -812 ne
rect 24829 -1148 24895 -812
rect 24829 -1204 24834 -1148
rect 24890 -1204 24895 -1148
rect 24829 -1228 24895 -1204
rect 24829 -1284 24834 -1228
rect 24890 -1284 24895 -1228
rect 24829 -1289 24895 -1284
rect 24963 -1148 25029 -572
rect 24963 -1204 24968 -1148
rect 25024 -1204 25029 -1148
rect 24963 -1228 25029 -1204
rect 24963 -1284 24968 -1228
rect 25024 -1284 25029 -1228
rect 24963 -1289 25029 -1284
rect 25089 -1316 25155 -211
rect 25089 -1372 25094 -1316
rect 25150 -1372 25155 -1316
rect 25089 -1396 25155 -1372
rect 25089 -1452 25094 -1396
rect 25150 -1452 25155 -1396
rect 25089 -1457 25155 -1452
rect 4845 -1913 4911 -1908
rect 4845 -1969 4850 -1913
rect 4906 -1969 4911 -1913
rect 4845 -1993 4911 -1969
rect 4845 -2049 4850 -1993
rect 4906 -2049 4911 -1993
rect 4845 -3715 4911 -2049
rect 4845 -3771 4850 -3715
rect 4906 -3771 4911 -3715
rect 4845 -3795 4911 -3771
rect 4845 -3851 4850 -3795
rect 4906 -3851 4911 -3795
rect 4845 -3860 4911 -3851
use sky130_fd_io__gpio_ovtv2_ctl_hld_i2c_fix  sky130_fd_io__gpio_ovtv2_ctl_hld_i2c_fix_0
timestamp 1683767628
transform -1 0 6601 0 1 10
box -165 -3 6151 2077
use sky130_fd_io__gpio_ovtv2_ctl_lsbank_i2c_fix  sky130_fd_io__gpio_ovtv2_ctl_lsbank_i2c_fix_0
timestamp 1683767628
transform 1 0 6541 0 1 72
box -6326 -939 21038 2015
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1683767628
transform -1 0 572 0 -1 2079
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_1
timestamp 1683767628
transform 1 0 1160 0 1 -2
box 107 226 240 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1683767628
transform -1 0 1034 0 -1 2079
box 107 226 460 873
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_0
timestamp 1683767628
transform 1 0 24705 0 -1 -811
box 107 226 460 873
<< labels >>
flabel metal2 s 26950 95 26988 181 3 FreeSans 200 0 0 0 DM_H[0]
port 2 nsew
flabel metal2 s 23713 91 23747 182 3 FreeSans 200 0 0 0 DM_H[1]
port 3 nsew
flabel metal2 s 22801 102 22844 196 3 FreeSans 200 0 0 0 DM_H[2]
port 4 nsew
flabel metal2 s 26656 96 26693 214 3 FreeSans 200 0 0 0 DM_H_N[0]
port 5 nsew
flabel metal2 s 24016 96 24046 224 3 FreeSans 200 0 0 0 DM_H_N[1]
port 6 nsew
flabel metal2 s 22513 90 22546 213 3 FreeSans 200 0 0 0 DM_H_N[2]
port 7 nsew
flabel metal2 s 25417 92 25454 199 3 FreeSans 200 0 0 0 DM[0]
port 8 nsew
flabel metal2 s 25248 88 25283 211 3 FreeSans 200 0 0 0 DM[1]
port 9 nsew
flabel metal2 s 21268 85 21309 177 3 FreeSans 200 0 0 0 DM[2]
port 10 nsew
flabel metal2 s 21101 81 21141 161 3 FreeSans 200 0 0 0 INP_DIS
port 11 nsew
flabel metal2 s 19865 85 19904 175 3 FreeSans 200 0 0 0 INP_DIS_H_N
port 12 nsew
flabel metal2 s 18654 84 18696 176 3 FreeSans 200 0 0 0 VTRIP_SEL_H
port 13 nsew
flabel metal2 s 17122 80 17161 165 3 FreeSans 200 0 0 0 VTRIP_SEL
port 14 nsew
flabel metal2 s 16956 83 16993 175 3 FreeSans 200 180 0 0 IB_MODE_SEL[0]
port 15 nsew
flabel metal2 s 12978 86 13016 180 3 FreeSans 200 0 0 0 IB_MODE_SEL[1]
port 16 nsew
flabel metal2 s 15421 84 15459 169 3 FreeSans 200 0 0 0 IB_MODE_SEL_H[0]
port 17 nsew
flabel metal2 s 14512 88 14550 198 3 FreeSans 200 0 0 0 IB_MODE_SEL_H[1]
port 18 nsew
flabel metal2 s 15720 91 15758 187 3 FreeSans 200 0 0 0 IB_MODE_SEL_H_N[0]
port 19 nsew
flabel metal2 s 14216 91 14252 218 3 FreeSans 200 0 0 0 IB_MODE_SEL_H_N[1]
port 20 nsew
flabel metal2 s 12817 94 12848 165 3 FreeSans 200 0 0 0 SLEW_CTL[0]
port 21 nsew
flabel metal2 s 8833 92 8868 185 3 FreeSans 200 0 0 0 SLEW_CTL[1]
port 22 nsew
flabel metal2 s 11274 82 11312 192 3 FreeSans 200 0 0 0 SLEW_CTL_H[0]
port 23 nsew
flabel metal2 s 10366 88 10404 197 3 FreeSans 200 0 0 0 SLEW_CTL_H[1]
port 24 nsew
flabel metal2 s 11572 89 11608 219 3 FreeSans 200 0 0 0 SLEW_CTL_H_N[0]
port 25 nsew
flabel metal2 s 10071 90 10110 227 3 FreeSans 200 0 0 0 SLEW_CTL_H_N[1]
port 26 nsew
flabel metal2 s 8662 86 8707 178 3 FreeSans 200 0 0 0 HYST_TRIM
port 27 nsew
flabel metal2 s 7128 79 7170 193 3 FreeSans 200 0 0 0 HYST_TRIM_H
port 28 nsew
flabel metal2 s 7423 78 7468 196 3 FreeSans 200 0 0 0 HYST_TRIM_H_N
port 29 nsew
flabel metal2 s 1069 6 1114 92 3 FreeSans 200 0 0 0 ENABLE_INP_H
port 30 nsew
flabel metal2 s 5061 5 5103 70 3 FreeSans 200 0 0 0 HLD_OVR
port 31 nsew
flabel metal1 s 1333 -54 1502 -13 3 FreeSans 200 0 0 0 HLD_I_H_N
port 33 nsew
flabel metal1 s 2321 1490 2442 1561 3 FreeSans 520 0 0 0 ENABLE_H
port 34 nsew
flabel metal1 s 1143 357 1282 393 3 FreeSans 200 0 0 0 OD_I_H_N
port 35 nsew
flabel metal1 s 10997 211 11468 379 3 FreeSans 200 0 0 0 VDDIO_Q
port 36 nsew
flabel metal1 s 11109 1913 11446 2058 3 FreeSans 200 0 0 0 VCCD
port 37 nsew
flabel metal1 s 11163 1208 11555 1356 3 FreeSans 200 0 0 0 VSSD
port 38 nsew
flabel metal1 s 25062 -950 25062 -950 0 FreeSans 440 0 0 0 VSSD
flabel metal1 s 24952 -1743 24952 -1743 0 FreeSans 440 0 0 0 VDDIO_Q
flabel metal1 s 3897 1427 3939 1510 3 FreeSans 520 0 0 0 HLD_I_OVR_H
port 39 nsew
flabel metal1 s 2357 1658 2379 1721 3 FreeSans 520 0 0 0 HLD_H_N
port 40 nsew
flabel metal1 s 24871 -1199 24871 -1199 0 FreeSans 440 90 0 0 ENABLE_INP_H
<< properties >>
string GDS_END 35939100
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 35909242
<< end >>
