magic
tech sky130A
magscale 1 2
timestamp 1683767628
use sky130_fd_pr__dfl1sd2__example_55959141808521  sky130_fd_pr__dfl1sd2__example_55959141808521_0
timestamp 1683767628
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808521  sky130_fd_pr__dfl1sd2__example_55959141808521_1
timestamp 1683767628
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808520  sky130_fd_pr__dfl1sd__example_55959141808520_0
timestamp 1683767628
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808520  sky130_fd_pr__dfl1sd__example_55959141808520_1
timestamp 1683767628
transform 1 0 412 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 47728748
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 47726794
<< end >>
