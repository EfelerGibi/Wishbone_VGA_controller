magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -47 769 4217 1263
<< mvpmos >>
rect 19 1044 2019 1144
rect 2151 1044 4151 1144
rect 19 888 2019 988
rect 2151 888 4151 988
<< mvpdiff >>
rect 19 1189 2019 1197
rect 19 1155 69 1189
rect 103 1155 137 1189
rect 171 1155 205 1189
rect 239 1155 273 1189
rect 307 1155 341 1189
rect 375 1155 409 1189
rect 443 1155 477 1189
rect 511 1155 545 1189
rect 579 1155 613 1189
rect 647 1155 681 1189
rect 715 1155 749 1189
rect 783 1155 817 1189
rect 851 1155 885 1189
rect 919 1155 953 1189
rect 987 1155 1021 1189
rect 1055 1155 1089 1189
rect 1123 1155 1157 1189
rect 1191 1155 1225 1189
rect 1259 1155 1293 1189
rect 1327 1155 1361 1189
rect 1395 1155 1429 1189
rect 1463 1155 1497 1189
rect 1531 1155 1565 1189
rect 1599 1155 1633 1189
rect 1667 1155 1701 1189
rect 1735 1155 1769 1189
rect 1803 1155 1837 1189
rect 1871 1155 1905 1189
rect 1939 1155 1973 1189
rect 2007 1155 2019 1189
rect 19 1144 2019 1155
rect 2151 1189 4151 1197
rect 2151 1155 2163 1189
rect 2197 1155 2231 1189
rect 2265 1155 2299 1189
rect 2333 1155 2367 1189
rect 2401 1155 2435 1189
rect 2469 1155 2503 1189
rect 2537 1155 2571 1189
rect 2605 1155 2639 1189
rect 2673 1155 2707 1189
rect 2741 1155 2775 1189
rect 2809 1155 2843 1189
rect 2877 1155 2911 1189
rect 2945 1155 2979 1189
rect 3013 1155 3047 1189
rect 3081 1155 3115 1189
rect 3149 1155 3183 1189
rect 3217 1155 3251 1189
rect 3285 1155 3319 1189
rect 3353 1155 3387 1189
rect 3421 1155 3455 1189
rect 3489 1155 3523 1189
rect 3557 1155 3591 1189
rect 3625 1155 3659 1189
rect 3693 1155 3727 1189
rect 3761 1155 3795 1189
rect 3829 1155 3863 1189
rect 3897 1155 3931 1189
rect 3965 1155 3999 1189
rect 4033 1155 4067 1189
rect 4101 1155 4151 1189
rect 2151 1144 4151 1155
rect 19 1033 2019 1044
rect 19 999 69 1033
rect 103 999 137 1033
rect 171 999 205 1033
rect 239 999 273 1033
rect 307 999 341 1033
rect 375 999 409 1033
rect 443 999 477 1033
rect 511 999 545 1033
rect 579 999 613 1033
rect 647 999 681 1033
rect 715 999 749 1033
rect 783 999 817 1033
rect 851 999 885 1033
rect 919 999 953 1033
rect 987 999 1021 1033
rect 1055 999 1089 1033
rect 1123 999 1157 1033
rect 1191 999 1225 1033
rect 1259 999 1293 1033
rect 1327 999 1361 1033
rect 1395 999 1429 1033
rect 1463 999 1497 1033
rect 1531 999 1565 1033
rect 1599 999 1633 1033
rect 1667 999 1701 1033
rect 1735 999 1769 1033
rect 1803 999 1837 1033
rect 1871 999 1905 1033
rect 1939 999 1973 1033
rect 2007 999 2019 1033
rect 19 988 2019 999
rect 2151 1033 4151 1044
rect 2151 999 2163 1033
rect 2197 999 2231 1033
rect 2265 999 2299 1033
rect 2333 999 2367 1033
rect 2401 999 2435 1033
rect 2469 999 2503 1033
rect 2537 999 2571 1033
rect 2605 999 2639 1033
rect 2673 999 2707 1033
rect 2741 999 2775 1033
rect 2809 999 2843 1033
rect 2877 999 2911 1033
rect 2945 999 2979 1033
rect 3013 999 3047 1033
rect 3081 999 3115 1033
rect 3149 999 3183 1033
rect 3217 999 3251 1033
rect 3285 999 3319 1033
rect 3353 999 3387 1033
rect 3421 999 3455 1033
rect 3489 999 3523 1033
rect 3557 999 3591 1033
rect 3625 999 3659 1033
rect 3693 999 3727 1033
rect 3761 999 3795 1033
rect 3829 999 3863 1033
rect 3897 999 3931 1033
rect 3965 999 3999 1033
rect 4033 999 4067 1033
rect 4101 999 4151 1033
rect 2151 988 4151 999
rect 19 877 2019 888
rect 19 843 69 877
rect 103 843 137 877
rect 171 843 205 877
rect 239 843 273 877
rect 307 843 341 877
rect 375 843 409 877
rect 443 843 477 877
rect 511 843 545 877
rect 579 843 613 877
rect 647 843 681 877
rect 715 843 749 877
rect 783 843 817 877
rect 851 843 885 877
rect 919 843 953 877
rect 987 843 1021 877
rect 1055 843 1089 877
rect 1123 843 1157 877
rect 1191 843 1225 877
rect 1259 843 1293 877
rect 1327 843 1361 877
rect 1395 843 1429 877
rect 1463 843 1497 877
rect 1531 843 1565 877
rect 1599 843 1633 877
rect 1667 843 1701 877
rect 1735 843 1769 877
rect 1803 843 1837 877
rect 1871 843 1905 877
rect 1939 843 1973 877
rect 2007 843 2019 877
rect 19 835 2019 843
rect 2151 877 4151 888
rect 2151 843 2163 877
rect 2197 843 2231 877
rect 2265 843 2299 877
rect 2333 843 2367 877
rect 2401 843 2435 877
rect 2469 843 2503 877
rect 2537 843 2571 877
rect 2605 843 2639 877
rect 2673 843 2707 877
rect 2741 843 2775 877
rect 2809 843 2843 877
rect 2877 843 2911 877
rect 2945 843 2979 877
rect 3013 843 3047 877
rect 3081 843 3115 877
rect 3149 843 3183 877
rect 3217 843 3251 877
rect 3285 843 3319 877
rect 3353 843 3387 877
rect 3421 843 3455 877
rect 3489 843 3523 877
rect 3557 843 3591 877
rect 3625 843 3659 877
rect 3693 843 3727 877
rect 3761 843 3795 877
rect 3829 843 3863 877
rect 3897 843 3931 877
rect 3965 843 3999 877
rect 4033 843 4067 877
rect 4101 843 4151 877
rect 2151 835 4151 843
<< mvpdiffc >>
rect 69 1155 103 1189
rect 137 1155 171 1189
rect 205 1155 239 1189
rect 273 1155 307 1189
rect 341 1155 375 1189
rect 409 1155 443 1189
rect 477 1155 511 1189
rect 545 1155 579 1189
rect 613 1155 647 1189
rect 681 1155 715 1189
rect 749 1155 783 1189
rect 817 1155 851 1189
rect 885 1155 919 1189
rect 953 1155 987 1189
rect 1021 1155 1055 1189
rect 1089 1155 1123 1189
rect 1157 1155 1191 1189
rect 1225 1155 1259 1189
rect 1293 1155 1327 1189
rect 1361 1155 1395 1189
rect 1429 1155 1463 1189
rect 1497 1155 1531 1189
rect 1565 1155 1599 1189
rect 1633 1155 1667 1189
rect 1701 1155 1735 1189
rect 1769 1155 1803 1189
rect 1837 1155 1871 1189
rect 1905 1155 1939 1189
rect 1973 1155 2007 1189
rect 2163 1155 2197 1189
rect 2231 1155 2265 1189
rect 2299 1155 2333 1189
rect 2367 1155 2401 1189
rect 2435 1155 2469 1189
rect 2503 1155 2537 1189
rect 2571 1155 2605 1189
rect 2639 1155 2673 1189
rect 2707 1155 2741 1189
rect 2775 1155 2809 1189
rect 2843 1155 2877 1189
rect 2911 1155 2945 1189
rect 2979 1155 3013 1189
rect 3047 1155 3081 1189
rect 3115 1155 3149 1189
rect 3183 1155 3217 1189
rect 3251 1155 3285 1189
rect 3319 1155 3353 1189
rect 3387 1155 3421 1189
rect 3455 1155 3489 1189
rect 3523 1155 3557 1189
rect 3591 1155 3625 1189
rect 3659 1155 3693 1189
rect 3727 1155 3761 1189
rect 3795 1155 3829 1189
rect 3863 1155 3897 1189
rect 3931 1155 3965 1189
rect 3999 1155 4033 1189
rect 4067 1155 4101 1189
rect 69 999 103 1033
rect 137 999 171 1033
rect 205 999 239 1033
rect 273 999 307 1033
rect 341 999 375 1033
rect 409 999 443 1033
rect 477 999 511 1033
rect 545 999 579 1033
rect 613 999 647 1033
rect 681 999 715 1033
rect 749 999 783 1033
rect 817 999 851 1033
rect 885 999 919 1033
rect 953 999 987 1033
rect 1021 999 1055 1033
rect 1089 999 1123 1033
rect 1157 999 1191 1033
rect 1225 999 1259 1033
rect 1293 999 1327 1033
rect 1361 999 1395 1033
rect 1429 999 1463 1033
rect 1497 999 1531 1033
rect 1565 999 1599 1033
rect 1633 999 1667 1033
rect 1701 999 1735 1033
rect 1769 999 1803 1033
rect 1837 999 1871 1033
rect 1905 999 1939 1033
rect 1973 999 2007 1033
rect 2163 999 2197 1033
rect 2231 999 2265 1033
rect 2299 999 2333 1033
rect 2367 999 2401 1033
rect 2435 999 2469 1033
rect 2503 999 2537 1033
rect 2571 999 2605 1033
rect 2639 999 2673 1033
rect 2707 999 2741 1033
rect 2775 999 2809 1033
rect 2843 999 2877 1033
rect 2911 999 2945 1033
rect 2979 999 3013 1033
rect 3047 999 3081 1033
rect 3115 999 3149 1033
rect 3183 999 3217 1033
rect 3251 999 3285 1033
rect 3319 999 3353 1033
rect 3387 999 3421 1033
rect 3455 999 3489 1033
rect 3523 999 3557 1033
rect 3591 999 3625 1033
rect 3659 999 3693 1033
rect 3727 999 3761 1033
rect 3795 999 3829 1033
rect 3863 999 3897 1033
rect 3931 999 3965 1033
rect 3999 999 4033 1033
rect 4067 999 4101 1033
rect 69 843 103 877
rect 137 843 171 877
rect 205 843 239 877
rect 273 843 307 877
rect 341 843 375 877
rect 409 843 443 877
rect 477 843 511 877
rect 545 843 579 877
rect 613 843 647 877
rect 681 843 715 877
rect 749 843 783 877
rect 817 843 851 877
rect 885 843 919 877
rect 953 843 987 877
rect 1021 843 1055 877
rect 1089 843 1123 877
rect 1157 843 1191 877
rect 1225 843 1259 877
rect 1293 843 1327 877
rect 1361 843 1395 877
rect 1429 843 1463 877
rect 1497 843 1531 877
rect 1565 843 1599 877
rect 1633 843 1667 877
rect 1701 843 1735 877
rect 1769 843 1803 877
rect 1837 843 1871 877
rect 1905 843 1939 877
rect 1973 843 2007 877
rect 2163 843 2197 877
rect 2231 843 2265 877
rect 2299 843 2333 877
rect 2367 843 2401 877
rect 2435 843 2469 877
rect 2503 843 2537 877
rect 2571 843 2605 877
rect 2639 843 2673 877
rect 2707 843 2741 877
rect 2775 843 2809 877
rect 2843 843 2877 877
rect 2911 843 2945 877
rect 2979 843 3013 877
rect 3047 843 3081 877
rect 3115 843 3149 877
rect 3183 843 3217 877
rect 3251 843 3285 877
rect 3319 843 3353 877
rect 3387 843 3421 877
rect 3455 843 3489 877
rect 3523 843 3557 877
rect 3591 843 3625 877
rect 3659 843 3693 877
rect 3727 843 3761 877
rect 3795 843 3829 877
rect 3863 843 3897 877
rect 3931 843 3965 877
rect 3999 843 4033 877
rect 4067 843 4101 877
<< poly >>
rect -80 1128 19 1144
rect -80 1094 -64 1128
rect -30 1094 19 1128
rect -80 1044 19 1094
rect 2019 1128 2151 1144
rect 2019 1094 2068 1128
rect 2102 1094 2151 1128
rect 2019 1044 2151 1094
rect 4151 1128 4257 1144
rect 4151 1094 4200 1128
rect 4234 1094 4257 1128
rect 4151 1044 4257 1094
rect -80 1033 0 1044
rect -80 999 -64 1033
rect -30 999 0 1033
rect -80 988 0 999
rect 2052 1033 2118 1044
rect 2052 999 2068 1033
rect 2102 999 2118 1033
rect 2052 988 2118 999
rect 4177 1033 4257 1044
rect 4177 999 4200 1033
rect 4234 999 4257 1033
rect 4177 988 4257 999
rect -80 938 19 988
rect -80 904 -64 938
rect -30 904 19 938
rect -80 888 19 904
rect 2019 938 2151 988
rect 2019 904 2068 938
rect 2102 904 2151 938
rect 2019 888 2151 904
rect 4151 938 4257 988
rect 4151 904 4200 938
rect 4234 904 4257 938
rect 4151 888 4257 904
<< polycont >>
rect -64 1094 -30 1128
rect 2068 1094 2102 1128
rect 4200 1094 4234 1128
rect -64 999 -30 1033
rect 2068 999 2102 1033
rect 4200 999 4234 1033
rect -64 904 -30 938
rect 2068 904 2102 938
rect 4200 904 4234 938
<< locali >>
rect 103 1155 117 1189
rect 171 1155 189 1189
rect 239 1155 261 1189
rect 307 1155 333 1189
rect 375 1155 405 1189
rect 443 1155 477 1189
rect 511 1155 545 1189
rect 583 1155 613 1189
rect 655 1155 681 1189
rect 727 1155 749 1189
rect 799 1155 817 1189
rect 871 1155 885 1189
rect 943 1155 953 1189
rect 1015 1155 1021 1189
rect 1087 1155 1089 1189
rect 1123 1155 1125 1189
rect 1191 1155 1197 1189
rect 1259 1155 1269 1189
rect 1327 1155 1341 1189
rect 1395 1155 1413 1189
rect 1463 1155 1485 1189
rect 1531 1155 1557 1189
rect 1599 1155 1629 1189
rect 1667 1155 1701 1189
rect 1735 1155 1769 1189
rect 1807 1155 1837 1189
rect 1879 1155 1905 1189
rect 1951 1155 1973 1189
rect 2197 1155 2219 1189
rect 2265 1155 2291 1189
rect 2333 1155 2363 1189
rect 2401 1155 2435 1189
rect 2469 1155 2503 1189
rect 2541 1155 2571 1189
rect 2613 1155 2639 1189
rect 2685 1155 2707 1189
rect 2757 1155 2775 1189
rect 2829 1155 2843 1189
rect 2901 1155 2911 1189
rect 2973 1155 2979 1189
rect 3045 1155 3047 1189
rect 3081 1155 3083 1189
rect 3149 1155 3155 1189
rect 3217 1155 3227 1189
rect 3285 1155 3299 1189
rect 3353 1155 3371 1189
rect 3421 1155 3443 1189
rect 3489 1155 3515 1189
rect 3557 1155 3587 1189
rect 3625 1155 3659 1189
rect 3693 1155 3727 1189
rect 3765 1155 3795 1189
rect 3837 1155 3863 1189
rect 3909 1155 3931 1189
rect 3981 1155 3999 1189
rect 4053 1155 4067 1189
rect -64 1128 -30 1144
rect 2057 1128 2113 1145
rect 2057 1117 2068 1128
rect -30 1094 2068 1117
rect 2102 1117 2113 1128
rect 4200 1128 4234 1144
rect 2102 1094 4200 1117
rect -64 1071 4234 1094
rect -64 1033 -30 1071
rect 2057 1033 2113 1071
rect 4200 1033 4234 1071
rect 103 999 117 1033
rect 171 999 189 1033
rect 239 999 261 1033
rect 307 999 333 1033
rect 375 999 405 1033
rect 443 999 477 1033
rect 511 999 545 1033
rect 583 999 613 1033
rect 655 999 681 1033
rect 727 999 749 1033
rect 799 999 817 1033
rect 871 999 885 1033
rect 943 999 953 1033
rect 1015 999 1021 1033
rect 1087 999 1089 1033
rect 1123 999 1125 1033
rect 1191 999 1197 1033
rect 1259 999 1269 1033
rect 1327 999 1341 1033
rect 1395 999 1413 1033
rect 1463 999 1485 1033
rect 1531 999 1557 1033
rect 1599 999 1629 1033
rect 1667 999 1701 1033
rect 1735 999 1769 1033
rect 1807 999 1837 1033
rect 1879 999 1905 1033
rect 1951 999 1973 1033
rect 2057 999 2068 1033
rect 2102 999 2113 1033
rect 2197 999 2219 1033
rect 2265 999 2291 1033
rect 2333 999 2363 1033
rect 2401 999 2435 1033
rect 2469 999 2503 1033
rect 2541 999 2571 1033
rect 2613 999 2639 1033
rect 2685 999 2707 1033
rect 2757 999 2775 1033
rect 2829 999 2843 1033
rect 2901 999 2911 1033
rect 2973 999 2979 1033
rect 3045 999 3047 1033
rect 3081 999 3083 1033
rect 3149 999 3155 1033
rect 3217 999 3227 1033
rect 3285 999 3299 1033
rect 3353 999 3371 1033
rect 3421 999 3443 1033
rect 3489 999 3515 1033
rect 3557 999 3587 1033
rect 3625 999 3659 1033
rect 3693 999 3727 1033
rect 3765 999 3795 1033
rect 3837 999 3863 1033
rect 3909 999 3931 1033
rect 3981 999 3999 1033
rect 4053 999 4067 1033
rect -64 961 -30 999
rect 2057 961 2113 999
rect 4200 961 4234 999
rect -64 955 4234 961
rect -64 938 2033 955
rect -30 921 2033 938
rect 2067 938 2105 955
rect 2067 921 2068 938
rect -30 915 2068 921
rect -64 888 -30 904
rect 2057 904 2068 915
rect 2102 921 2105 938
rect 2139 938 4234 955
rect 2139 921 4200 938
rect 2102 915 4200 921
rect 2102 904 2113 915
rect 2057 888 2113 904
rect 4200 888 4234 904
rect 103 843 117 877
rect 171 843 189 877
rect 239 843 261 877
rect 307 843 333 877
rect 375 843 405 877
rect 443 843 477 877
rect 511 843 545 877
rect 583 843 613 877
rect 655 843 681 877
rect 727 843 749 877
rect 799 843 817 877
rect 871 843 885 877
rect 943 843 953 877
rect 1015 843 1021 877
rect 1087 843 1089 877
rect 1123 843 1125 877
rect 1191 843 1197 877
rect 1259 843 1269 877
rect 1327 843 1341 877
rect 1395 843 1413 877
rect 1463 843 1485 877
rect 1531 843 1557 877
rect 1599 843 1629 877
rect 1667 843 1701 877
rect 1735 843 1769 877
rect 1807 843 1837 877
rect 1879 843 1905 877
rect 1951 843 1973 877
rect 2197 843 2219 877
rect 2265 843 2291 877
rect 2333 843 2363 877
rect 2401 843 2435 877
rect 2469 843 2503 877
rect 2541 843 2571 877
rect 2613 843 2639 877
rect 2685 843 2707 877
rect 2757 843 2775 877
rect 2829 843 2843 877
rect 2901 843 2911 877
rect 2973 843 2979 877
rect 3045 843 3047 877
rect 3081 843 3083 877
rect 3149 843 3155 877
rect 3217 843 3227 877
rect 3285 843 3299 877
rect 3353 843 3371 877
rect 3421 843 3443 877
rect 3489 843 3515 877
rect 3557 843 3587 877
rect 3625 843 3659 877
rect 3693 843 3727 877
rect 3765 843 3795 877
rect 3837 843 3863 877
rect 3909 843 3931 877
rect 3981 843 3999 877
rect 4053 843 4067 877
<< viali >>
rect 45 1155 69 1189
rect 69 1155 79 1189
rect 117 1155 137 1189
rect 137 1155 151 1189
rect 189 1155 205 1189
rect 205 1155 223 1189
rect 261 1155 273 1189
rect 273 1155 295 1189
rect 333 1155 341 1189
rect 341 1155 367 1189
rect 405 1155 409 1189
rect 409 1155 439 1189
rect 477 1155 511 1189
rect 549 1155 579 1189
rect 579 1155 583 1189
rect 621 1155 647 1189
rect 647 1155 655 1189
rect 693 1155 715 1189
rect 715 1155 727 1189
rect 765 1155 783 1189
rect 783 1155 799 1189
rect 837 1155 851 1189
rect 851 1155 871 1189
rect 909 1155 919 1189
rect 919 1155 943 1189
rect 981 1155 987 1189
rect 987 1155 1015 1189
rect 1053 1155 1055 1189
rect 1055 1155 1087 1189
rect 1125 1155 1157 1189
rect 1157 1155 1159 1189
rect 1197 1155 1225 1189
rect 1225 1155 1231 1189
rect 1269 1155 1293 1189
rect 1293 1155 1303 1189
rect 1341 1155 1361 1189
rect 1361 1155 1375 1189
rect 1413 1155 1429 1189
rect 1429 1155 1447 1189
rect 1485 1155 1497 1189
rect 1497 1155 1519 1189
rect 1557 1155 1565 1189
rect 1565 1155 1591 1189
rect 1629 1155 1633 1189
rect 1633 1155 1663 1189
rect 1701 1155 1735 1189
rect 1773 1155 1803 1189
rect 1803 1155 1807 1189
rect 1845 1155 1871 1189
rect 1871 1155 1879 1189
rect 1917 1155 1939 1189
rect 1939 1155 1951 1189
rect 1989 1155 2007 1189
rect 2007 1155 2023 1189
rect 2147 1155 2163 1189
rect 2163 1155 2181 1189
rect 2219 1155 2231 1189
rect 2231 1155 2253 1189
rect 2291 1155 2299 1189
rect 2299 1155 2325 1189
rect 2363 1155 2367 1189
rect 2367 1155 2397 1189
rect 2435 1155 2469 1189
rect 2507 1155 2537 1189
rect 2537 1155 2541 1189
rect 2579 1155 2605 1189
rect 2605 1155 2613 1189
rect 2651 1155 2673 1189
rect 2673 1155 2685 1189
rect 2723 1155 2741 1189
rect 2741 1155 2757 1189
rect 2795 1155 2809 1189
rect 2809 1155 2829 1189
rect 2867 1155 2877 1189
rect 2877 1155 2901 1189
rect 2939 1155 2945 1189
rect 2945 1155 2973 1189
rect 3011 1155 3013 1189
rect 3013 1155 3045 1189
rect 3083 1155 3115 1189
rect 3115 1155 3117 1189
rect 3155 1155 3183 1189
rect 3183 1155 3189 1189
rect 3227 1155 3251 1189
rect 3251 1155 3261 1189
rect 3299 1155 3319 1189
rect 3319 1155 3333 1189
rect 3371 1155 3387 1189
rect 3387 1155 3405 1189
rect 3443 1155 3455 1189
rect 3455 1155 3477 1189
rect 3515 1155 3523 1189
rect 3523 1155 3549 1189
rect 3587 1155 3591 1189
rect 3591 1155 3621 1189
rect 3659 1155 3693 1189
rect 3731 1155 3761 1189
rect 3761 1155 3765 1189
rect 3803 1155 3829 1189
rect 3829 1155 3837 1189
rect 3875 1155 3897 1189
rect 3897 1155 3909 1189
rect 3947 1155 3965 1189
rect 3965 1155 3981 1189
rect 4019 1155 4033 1189
rect 4033 1155 4053 1189
rect 4091 1155 4101 1189
rect 4101 1155 4125 1189
rect 45 999 69 1033
rect 69 999 79 1033
rect 117 999 137 1033
rect 137 999 151 1033
rect 189 999 205 1033
rect 205 999 223 1033
rect 261 999 273 1033
rect 273 999 295 1033
rect 333 999 341 1033
rect 341 999 367 1033
rect 405 999 409 1033
rect 409 999 439 1033
rect 477 999 511 1033
rect 549 999 579 1033
rect 579 999 583 1033
rect 621 999 647 1033
rect 647 999 655 1033
rect 693 999 715 1033
rect 715 999 727 1033
rect 765 999 783 1033
rect 783 999 799 1033
rect 837 999 851 1033
rect 851 999 871 1033
rect 909 999 919 1033
rect 919 999 943 1033
rect 981 999 987 1033
rect 987 999 1015 1033
rect 1053 999 1055 1033
rect 1055 999 1087 1033
rect 1125 999 1157 1033
rect 1157 999 1159 1033
rect 1197 999 1225 1033
rect 1225 999 1231 1033
rect 1269 999 1293 1033
rect 1293 999 1303 1033
rect 1341 999 1361 1033
rect 1361 999 1375 1033
rect 1413 999 1429 1033
rect 1429 999 1447 1033
rect 1485 999 1497 1033
rect 1497 999 1519 1033
rect 1557 999 1565 1033
rect 1565 999 1591 1033
rect 1629 999 1633 1033
rect 1633 999 1663 1033
rect 1701 999 1735 1033
rect 1773 999 1803 1033
rect 1803 999 1807 1033
rect 1845 999 1871 1033
rect 1871 999 1879 1033
rect 1917 999 1939 1033
rect 1939 999 1951 1033
rect 1989 999 2007 1033
rect 2007 999 2023 1033
rect 2147 999 2163 1033
rect 2163 999 2181 1033
rect 2219 999 2231 1033
rect 2231 999 2253 1033
rect 2291 999 2299 1033
rect 2299 999 2325 1033
rect 2363 999 2367 1033
rect 2367 999 2397 1033
rect 2435 999 2469 1033
rect 2507 999 2537 1033
rect 2537 999 2541 1033
rect 2579 999 2605 1033
rect 2605 999 2613 1033
rect 2651 999 2673 1033
rect 2673 999 2685 1033
rect 2723 999 2741 1033
rect 2741 999 2757 1033
rect 2795 999 2809 1033
rect 2809 999 2829 1033
rect 2867 999 2877 1033
rect 2877 999 2901 1033
rect 2939 999 2945 1033
rect 2945 999 2973 1033
rect 3011 999 3013 1033
rect 3013 999 3045 1033
rect 3083 999 3115 1033
rect 3115 999 3117 1033
rect 3155 999 3183 1033
rect 3183 999 3189 1033
rect 3227 999 3251 1033
rect 3251 999 3261 1033
rect 3299 999 3319 1033
rect 3319 999 3333 1033
rect 3371 999 3387 1033
rect 3387 999 3405 1033
rect 3443 999 3455 1033
rect 3455 999 3477 1033
rect 3515 999 3523 1033
rect 3523 999 3549 1033
rect 3587 999 3591 1033
rect 3591 999 3621 1033
rect 3659 999 3693 1033
rect 3731 999 3761 1033
rect 3761 999 3765 1033
rect 3803 999 3829 1033
rect 3829 999 3837 1033
rect 3875 999 3897 1033
rect 3897 999 3909 1033
rect 3947 999 3965 1033
rect 3965 999 3981 1033
rect 4019 999 4033 1033
rect 4033 999 4053 1033
rect 4091 999 4101 1033
rect 4101 999 4125 1033
rect 2033 921 2067 955
rect 2105 921 2139 955
rect 45 843 69 877
rect 69 843 79 877
rect 117 843 137 877
rect 137 843 151 877
rect 189 843 205 877
rect 205 843 223 877
rect 261 843 273 877
rect 273 843 295 877
rect 333 843 341 877
rect 341 843 367 877
rect 405 843 409 877
rect 409 843 439 877
rect 477 843 511 877
rect 549 843 579 877
rect 579 843 583 877
rect 621 843 647 877
rect 647 843 655 877
rect 693 843 715 877
rect 715 843 727 877
rect 765 843 783 877
rect 783 843 799 877
rect 837 843 851 877
rect 851 843 871 877
rect 909 843 919 877
rect 919 843 943 877
rect 981 843 987 877
rect 987 843 1015 877
rect 1053 843 1055 877
rect 1055 843 1087 877
rect 1125 843 1157 877
rect 1157 843 1159 877
rect 1197 843 1225 877
rect 1225 843 1231 877
rect 1269 843 1293 877
rect 1293 843 1303 877
rect 1341 843 1361 877
rect 1361 843 1375 877
rect 1413 843 1429 877
rect 1429 843 1447 877
rect 1485 843 1497 877
rect 1497 843 1519 877
rect 1557 843 1565 877
rect 1565 843 1591 877
rect 1629 843 1633 877
rect 1633 843 1663 877
rect 1701 843 1735 877
rect 1773 843 1803 877
rect 1803 843 1807 877
rect 1845 843 1871 877
rect 1871 843 1879 877
rect 1917 843 1939 877
rect 1939 843 1951 877
rect 1989 843 2007 877
rect 2007 843 2023 877
rect 2147 843 2163 877
rect 2163 843 2181 877
rect 2219 843 2231 877
rect 2231 843 2253 877
rect 2291 843 2299 877
rect 2299 843 2325 877
rect 2363 843 2367 877
rect 2367 843 2397 877
rect 2435 843 2469 877
rect 2507 843 2537 877
rect 2537 843 2541 877
rect 2579 843 2605 877
rect 2605 843 2613 877
rect 2651 843 2673 877
rect 2673 843 2685 877
rect 2723 843 2741 877
rect 2741 843 2757 877
rect 2795 843 2809 877
rect 2809 843 2829 877
rect 2867 843 2877 877
rect 2877 843 2901 877
rect 2939 843 2945 877
rect 2945 843 2973 877
rect 3011 843 3013 877
rect 3013 843 3045 877
rect 3083 843 3115 877
rect 3115 843 3117 877
rect 3155 843 3183 877
rect 3183 843 3189 877
rect 3227 843 3251 877
rect 3251 843 3261 877
rect 3299 843 3319 877
rect 3319 843 3333 877
rect 3371 843 3387 877
rect 3387 843 3405 877
rect 3443 843 3455 877
rect 3455 843 3477 877
rect 3515 843 3523 877
rect 3523 843 3549 877
rect 3587 843 3591 877
rect 3591 843 3621 877
rect 3659 843 3693 877
rect 3731 843 3761 877
rect 3761 843 3765 877
rect 3803 843 3829 877
rect 3829 843 3837 877
rect 3875 843 3897 877
rect 3897 843 3909 877
rect 3947 843 3965 877
rect 3965 843 3981 877
rect 4019 843 4033 877
rect 4033 843 4053 877
rect 4091 843 4101 877
rect 4101 843 4125 877
<< metal1 >>
rect 33 1190 4139 1214
rect 33 1138 41 1190
rect 93 1138 112 1190
rect 164 1138 183 1190
rect 235 1138 254 1190
rect 306 1138 325 1190
rect 377 1138 396 1190
rect 448 1138 466 1190
rect 518 1138 536 1190
rect 588 1138 606 1190
rect 658 1138 676 1190
rect 728 1189 3446 1190
rect 3498 1189 3516 1190
rect 728 1155 765 1189
rect 799 1155 837 1189
rect 871 1155 909 1189
rect 943 1155 981 1189
rect 1015 1155 1053 1189
rect 1087 1155 1125 1189
rect 1159 1155 1197 1189
rect 1231 1155 1269 1189
rect 1303 1155 1341 1189
rect 1375 1155 1413 1189
rect 1447 1155 1485 1189
rect 1519 1155 1557 1189
rect 1591 1155 1629 1189
rect 1663 1155 1701 1189
rect 1735 1155 1773 1189
rect 1807 1155 1845 1189
rect 1879 1155 1917 1189
rect 1951 1155 1989 1189
rect 2023 1155 2147 1189
rect 2181 1155 2219 1189
rect 2253 1155 2291 1189
rect 2325 1155 2363 1189
rect 2397 1155 2435 1189
rect 2469 1155 2507 1189
rect 2541 1155 2579 1189
rect 2613 1155 2651 1189
rect 2685 1155 2723 1189
rect 2757 1155 2795 1189
rect 2829 1155 2867 1189
rect 2901 1155 2939 1189
rect 2973 1155 3011 1189
rect 3045 1155 3083 1189
rect 3117 1155 3155 1189
rect 3189 1155 3227 1189
rect 3261 1155 3299 1189
rect 3333 1155 3371 1189
rect 3405 1155 3443 1189
rect 3498 1155 3515 1189
rect 728 1138 3446 1155
rect 3498 1138 3516 1155
rect 3568 1138 3586 1190
rect 3638 1138 3656 1190
rect 3708 1138 3726 1190
rect 3778 1138 3797 1190
rect 3849 1138 3868 1190
rect 3920 1138 3939 1190
rect 3991 1138 4010 1190
rect 4062 1138 4081 1190
rect 4133 1138 4139 1190
rect 33 1114 4139 1138
rect 834 1039 840 1042
rect 33 1033 840 1039
rect 33 999 45 1033
rect 79 999 117 1033
rect 151 999 189 1033
rect 223 999 261 1033
rect 295 999 333 1033
rect 367 999 405 1033
rect 439 999 477 1033
rect 511 999 549 1033
rect 583 999 621 1033
rect 655 999 693 1033
rect 727 999 765 1033
rect 799 999 837 1033
rect 33 993 840 999
rect 834 990 840 993
rect 892 990 908 1042
rect 960 990 976 1042
rect 1028 990 1044 1042
rect 1096 990 1112 1042
rect 1164 990 1180 1042
rect 1232 990 1247 1042
rect 1299 1033 1314 1042
rect 1366 1033 1381 1042
rect 1433 1033 1448 1042
rect 1500 1039 1506 1042
rect 2338 1039 2344 1042
rect 1500 1033 2035 1039
rect 1303 999 1314 1033
rect 1375 999 1381 1033
rect 1447 999 1448 1033
rect 1519 999 1557 1033
rect 1591 999 1629 1033
rect 1663 999 1701 1033
rect 1735 999 1773 1033
rect 1807 999 1845 1033
rect 1879 999 1917 1033
rect 1951 999 1989 1033
rect 2023 999 2035 1033
rect 1299 990 1314 999
rect 1366 990 1381 999
rect 1433 990 1448 999
rect 1500 993 2035 999
rect 2135 1033 2344 1039
rect 2396 1033 2414 1042
rect 2466 1033 2484 1042
rect 2536 1033 2554 1042
rect 2606 1033 2624 1042
rect 2676 1033 2695 1042
rect 2747 1039 2753 1042
rect 2747 1033 4137 1039
rect 2135 999 2147 1033
rect 2181 999 2219 1033
rect 2253 999 2291 1033
rect 2325 999 2344 1033
rect 2397 999 2414 1033
rect 2469 999 2484 1033
rect 2541 999 2554 1033
rect 2613 999 2624 1033
rect 2685 999 2695 1033
rect 2757 999 2795 1033
rect 2829 999 2867 1033
rect 2901 999 2939 1033
rect 2973 999 3011 1033
rect 3045 999 3083 1033
rect 3117 999 3155 1033
rect 3189 999 3227 1033
rect 3261 999 3299 1033
rect 3333 999 3371 1033
rect 3405 999 3443 1033
rect 3477 999 3515 1033
rect 3549 999 3587 1033
rect 3621 999 3659 1033
rect 3693 999 3731 1033
rect 3765 999 3803 1033
rect 3837 999 3875 1033
rect 3909 999 3947 1033
rect 3981 999 4019 1033
rect 4053 999 4091 1033
rect 4125 999 4137 1033
rect 2135 993 2344 999
rect 1500 990 1506 993
rect 2338 990 2344 993
rect 2396 990 2414 999
rect 2466 990 2484 999
rect 2536 990 2554 999
rect 2606 990 2624 999
rect 2676 990 2695 999
rect 2747 993 4137 999
rect 2747 990 2753 993
rect 33 894 1963 918
rect 33 842 41 894
rect 93 842 112 894
rect 164 842 183 894
rect 235 842 254 894
rect 306 842 325 894
rect 377 842 396 894
rect 448 842 466 894
rect 518 842 536 894
rect 588 842 606 894
rect 658 842 676 894
rect 728 883 1963 894
tri 1963 883 1998 918 sw
rect 2021 912 2027 964
rect 2079 912 2093 964
rect 2145 912 2151 964
tri 2240 912 2246 918 se
rect 2246 912 4262 918
tri 2211 883 2240 912 se
rect 2240 894 4262 912
rect 2240 883 3446 894
rect 728 877 3446 883
rect 3498 877 3516 894
rect 728 843 765 877
rect 799 843 837 877
rect 871 843 909 877
rect 943 843 981 877
rect 1015 843 1053 877
rect 1087 843 1125 877
rect 1159 843 1197 877
rect 1231 843 1269 877
rect 1303 843 1341 877
rect 1375 843 1413 877
rect 1447 843 1485 877
rect 1519 843 1557 877
rect 1591 843 1629 877
rect 1663 843 1701 877
rect 1735 843 1773 877
rect 1807 843 1845 877
rect 1879 843 1917 877
rect 1951 843 1989 877
rect 2023 843 2147 877
rect 2181 843 2219 877
rect 2253 843 2291 877
rect 2325 843 2363 877
rect 2397 843 2435 877
rect 2469 843 2507 877
rect 2541 843 2579 877
rect 2613 843 2651 877
rect 2685 843 2723 877
rect 2757 843 2795 877
rect 2829 843 2867 877
rect 2901 843 2939 877
rect 2973 843 3011 877
rect 3045 843 3083 877
rect 3117 843 3155 877
rect 3189 843 3227 877
rect 3261 843 3299 877
rect 3333 843 3371 877
rect 3405 843 3443 877
rect 3498 843 3515 877
rect 728 842 3446 843
rect 3498 842 3516 843
rect 3568 842 3586 894
rect 3638 842 3656 894
rect 3708 842 3726 894
rect 3778 842 3797 894
rect 3849 842 3868 894
rect 3920 842 3939 894
rect 3991 842 4010 894
rect 4062 842 4081 894
rect 4133 842 4262 894
rect 33 818 4262 842
<< via1 >>
rect 41 1189 93 1190
rect 41 1155 45 1189
rect 45 1155 79 1189
rect 79 1155 93 1189
rect 41 1138 93 1155
rect 112 1189 164 1190
rect 112 1155 117 1189
rect 117 1155 151 1189
rect 151 1155 164 1189
rect 112 1138 164 1155
rect 183 1189 235 1190
rect 183 1155 189 1189
rect 189 1155 223 1189
rect 223 1155 235 1189
rect 183 1138 235 1155
rect 254 1189 306 1190
rect 254 1155 261 1189
rect 261 1155 295 1189
rect 295 1155 306 1189
rect 254 1138 306 1155
rect 325 1189 377 1190
rect 325 1155 333 1189
rect 333 1155 367 1189
rect 367 1155 377 1189
rect 325 1138 377 1155
rect 396 1189 448 1190
rect 396 1155 405 1189
rect 405 1155 439 1189
rect 439 1155 448 1189
rect 396 1138 448 1155
rect 466 1189 518 1190
rect 466 1155 477 1189
rect 477 1155 511 1189
rect 511 1155 518 1189
rect 466 1138 518 1155
rect 536 1189 588 1190
rect 536 1155 549 1189
rect 549 1155 583 1189
rect 583 1155 588 1189
rect 536 1138 588 1155
rect 606 1189 658 1190
rect 606 1155 621 1189
rect 621 1155 655 1189
rect 655 1155 658 1189
rect 606 1138 658 1155
rect 676 1189 728 1190
rect 3446 1189 3498 1190
rect 3516 1189 3568 1190
rect 676 1155 693 1189
rect 693 1155 727 1189
rect 727 1155 728 1189
rect 3446 1155 3477 1189
rect 3477 1155 3498 1189
rect 3516 1155 3549 1189
rect 3549 1155 3568 1189
rect 676 1138 728 1155
rect 3446 1138 3498 1155
rect 3516 1138 3568 1155
rect 3586 1189 3638 1190
rect 3586 1155 3587 1189
rect 3587 1155 3621 1189
rect 3621 1155 3638 1189
rect 3586 1138 3638 1155
rect 3656 1189 3708 1190
rect 3656 1155 3659 1189
rect 3659 1155 3693 1189
rect 3693 1155 3708 1189
rect 3656 1138 3708 1155
rect 3726 1189 3778 1190
rect 3726 1155 3731 1189
rect 3731 1155 3765 1189
rect 3765 1155 3778 1189
rect 3726 1138 3778 1155
rect 3797 1189 3849 1190
rect 3797 1155 3803 1189
rect 3803 1155 3837 1189
rect 3837 1155 3849 1189
rect 3797 1138 3849 1155
rect 3868 1189 3920 1190
rect 3868 1155 3875 1189
rect 3875 1155 3909 1189
rect 3909 1155 3920 1189
rect 3868 1138 3920 1155
rect 3939 1189 3991 1190
rect 3939 1155 3947 1189
rect 3947 1155 3981 1189
rect 3981 1155 3991 1189
rect 3939 1138 3991 1155
rect 4010 1189 4062 1190
rect 4010 1155 4019 1189
rect 4019 1155 4053 1189
rect 4053 1155 4062 1189
rect 4010 1138 4062 1155
rect 4081 1189 4133 1190
rect 4081 1155 4091 1189
rect 4091 1155 4125 1189
rect 4125 1155 4133 1189
rect 4081 1138 4133 1155
rect 840 1033 892 1042
rect 840 999 871 1033
rect 871 999 892 1033
rect 840 990 892 999
rect 908 1033 960 1042
rect 908 999 909 1033
rect 909 999 943 1033
rect 943 999 960 1033
rect 908 990 960 999
rect 976 1033 1028 1042
rect 976 999 981 1033
rect 981 999 1015 1033
rect 1015 999 1028 1033
rect 976 990 1028 999
rect 1044 1033 1096 1042
rect 1044 999 1053 1033
rect 1053 999 1087 1033
rect 1087 999 1096 1033
rect 1044 990 1096 999
rect 1112 1033 1164 1042
rect 1112 999 1125 1033
rect 1125 999 1159 1033
rect 1159 999 1164 1033
rect 1112 990 1164 999
rect 1180 1033 1232 1042
rect 1180 999 1197 1033
rect 1197 999 1231 1033
rect 1231 999 1232 1033
rect 1180 990 1232 999
rect 1247 1033 1299 1042
rect 1314 1033 1366 1042
rect 1381 1033 1433 1042
rect 1448 1033 1500 1042
rect 1247 999 1269 1033
rect 1269 999 1299 1033
rect 1314 999 1341 1033
rect 1341 999 1366 1033
rect 1381 999 1413 1033
rect 1413 999 1433 1033
rect 1448 999 1485 1033
rect 1485 999 1500 1033
rect 1247 990 1299 999
rect 1314 990 1366 999
rect 1381 990 1433 999
rect 1448 990 1500 999
rect 2344 1033 2396 1042
rect 2414 1033 2466 1042
rect 2484 1033 2536 1042
rect 2554 1033 2606 1042
rect 2624 1033 2676 1042
rect 2695 1033 2747 1042
rect 2344 999 2363 1033
rect 2363 999 2396 1033
rect 2414 999 2435 1033
rect 2435 999 2466 1033
rect 2484 999 2507 1033
rect 2507 999 2536 1033
rect 2554 999 2579 1033
rect 2579 999 2606 1033
rect 2624 999 2651 1033
rect 2651 999 2676 1033
rect 2695 999 2723 1033
rect 2723 999 2747 1033
rect 2344 990 2396 999
rect 2414 990 2466 999
rect 2484 990 2536 999
rect 2554 990 2606 999
rect 2624 990 2676 999
rect 2695 990 2747 999
rect 41 877 93 894
rect 41 843 45 877
rect 45 843 79 877
rect 79 843 93 877
rect 41 842 93 843
rect 112 877 164 894
rect 112 843 117 877
rect 117 843 151 877
rect 151 843 164 877
rect 112 842 164 843
rect 183 877 235 894
rect 183 843 189 877
rect 189 843 223 877
rect 223 843 235 877
rect 183 842 235 843
rect 254 877 306 894
rect 254 843 261 877
rect 261 843 295 877
rect 295 843 306 877
rect 254 842 306 843
rect 325 877 377 894
rect 325 843 333 877
rect 333 843 367 877
rect 367 843 377 877
rect 325 842 377 843
rect 396 877 448 894
rect 396 843 405 877
rect 405 843 439 877
rect 439 843 448 877
rect 396 842 448 843
rect 466 877 518 894
rect 466 843 477 877
rect 477 843 511 877
rect 511 843 518 877
rect 466 842 518 843
rect 536 877 588 894
rect 536 843 549 877
rect 549 843 583 877
rect 583 843 588 877
rect 536 842 588 843
rect 606 877 658 894
rect 606 843 621 877
rect 621 843 655 877
rect 655 843 658 877
rect 606 842 658 843
rect 676 877 728 894
rect 2027 955 2079 964
rect 2027 921 2033 955
rect 2033 921 2067 955
rect 2067 921 2079 955
rect 2027 912 2079 921
rect 2093 955 2145 964
rect 2093 921 2105 955
rect 2105 921 2139 955
rect 2139 921 2145 955
rect 2093 912 2145 921
rect 3446 877 3498 894
rect 3516 877 3568 894
rect 676 843 693 877
rect 693 843 727 877
rect 727 843 728 877
rect 3446 843 3477 877
rect 3477 843 3498 877
rect 3516 843 3549 877
rect 3549 843 3568 877
rect 676 842 728 843
rect 3446 842 3498 843
rect 3516 842 3568 843
rect 3586 877 3638 894
rect 3586 843 3587 877
rect 3587 843 3621 877
rect 3621 843 3638 877
rect 3586 842 3638 843
rect 3656 877 3708 894
rect 3656 843 3659 877
rect 3659 843 3693 877
rect 3693 843 3708 877
rect 3656 842 3708 843
rect 3726 877 3778 894
rect 3726 843 3731 877
rect 3731 843 3765 877
rect 3765 843 3778 877
rect 3726 842 3778 843
rect 3797 877 3849 894
rect 3797 843 3803 877
rect 3803 843 3837 877
rect 3837 843 3849 877
rect 3797 842 3849 843
rect 3868 877 3920 894
rect 3868 843 3875 877
rect 3875 843 3909 877
rect 3909 843 3920 877
rect 3868 842 3920 843
rect 3939 877 3991 894
rect 3939 843 3947 877
rect 3947 843 3981 877
rect 3981 843 3991 877
rect 3939 842 3991 843
rect 4010 877 4062 894
rect 4010 843 4019 877
rect 4019 843 4053 877
rect 4053 843 4062 877
rect 4010 842 4062 843
rect 4081 877 4133 894
rect 4081 843 4091 877
rect 4091 843 4125 877
rect 4125 843 4133 877
rect 4081 842 4133 843
<< metal2 >>
rect 35 1190 734 1220
rect 35 1138 41 1190
rect 93 1138 112 1190
rect 164 1138 183 1190
rect 235 1138 254 1190
rect 306 1138 325 1190
rect 377 1138 396 1190
rect 448 1138 466 1190
rect 518 1138 536 1190
rect 588 1138 606 1190
rect 658 1138 676 1190
rect 728 1138 734 1190
rect 35 894 734 1138
rect 834 1042 1508 1220
rect 834 990 840 1042
rect 892 990 908 1042
rect 960 990 976 1042
rect 1028 990 1044 1042
rect 1096 990 1112 1042
rect 1164 990 1180 1042
rect 1232 990 1247 1042
rect 1299 990 1314 1042
rect 1366 990 1381 1042
rect 1433 990 1448 1042
rect 1500 990 1508 1042
rect 834 895 1508 990
rect 2021 964 2151 1214
rect 3440 1190 4139 1220
rect 3440 1138 3446 1190
rect 3498 1138 3516 1190
rect 3568 1138 3586 1190
rect 3638 1138 3656 1190
rect 3708 1138 3726 1190
rect 3778 1138 3797 1190
rect 3849 1138 3868 1190
rect 3920 1138 3939 1190
rect 3991 1138 4010 1190
rect 4062 1138 4081 1190
rect 4133 1138 4139 1190
rect 2021 912 2027 964
rect 2079 912 2093 964
rect 2145 912 2151 964
rect 35 842 41 894
rect 93 842 112 894
rect 164 842 183 894
rect 235 842 254 894
rect 306 842 325 894
rect 377 842 396 894
rect 448 842 466 894
rect 518 842 536 894
rect 588 842 606 894
rect 658 842 676 894
rect 728 842 734 894
rect 35 817 734 842
rect 2021 815 2151 912
rect 2336 1042 2753 1111
rect 2336 990 2344 1042
rect 2396 990 2414 1042
rect 2466 990 2484 1042
rect 2536 990 2554 1042
rect 2606 990 2624 1042
rect 2676 990 2695 1042
rect 2747 990 2753 1042
rect 2336 819 2753 990
rect 3440 894 4139 1138
rect 3440 842 3446 894
rect 3498 842 3516 894
rect 3568 842 3586 894
rect 3638 842 3656 894
rect 3708 842 3726 894
rect 3778 842 3797 894
rect 3849 842 3868 894
rect 3920 842 3939 894
rect 3991 842 4010 894
rect 4062 842 4081 894
rect 4133 842 4139 894
rect 3440 818 4139 842
use sky130_fd_pr__pfet_01v8__example_55959141808526  sky130_fd_pr__pfet_01v8__example_55959141808526_0
timestamp 1683767628
transform 0 1 2151 1 0 1044
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808526  sky130_fd_pr__pfet_01v8__example_55959141808526_1
timestamp 1683767628
transform 0 -1 2019 1 0 1044
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808526  sky130_fd_pr__pfet_01v8__example_55959141808526_2
timestamp 1683767628
transform 0 -1 2019 1 0 888
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808526  sky130_fd_pr__pfet_01v8__example_55959141808526_3
timestamp 1683767628
transform 0 1 2151 1 0 888
box -1 0 101 1
<< properties >>
string GDS_END 47717102
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 47709410
<< end >>
