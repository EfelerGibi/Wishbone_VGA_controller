magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 134 157 884 203
rect 37 21 884 157
rect 37 17 59 21
rect 25 -17 59 17
<< locali >>
rect 17 199 115 340
rect 816 299 903 493
rect 831 165 903 299
rect 816 51 903 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 17 408 105 493
rect 139 442 216 527
rect 17 374 216 408
rect 149 265 216 374
rect 250 335 304 493
rect 338 408 388 493
rect 422 442 499 527
rect 338 369 499 408
rect 250 299 395 335
rect 149 199 231 265
rect 265 199 395 299
rect 429 265 499 369
rect 533 335 583 493
rect 617 408 671 493
rect 705 442 782 527
rect 617 369 782 408
rect 533 299 678 335
rect 429 199 514 265
rect 548 199 678 299
rect 712 265 782 369
rect 712 199 797 265
rect 149 165 216 199
rect 265 165 304 199
rect 429 165 499 199
rect 548 165 583 199
rect 712 165 782 199
rect 17 131 216 165
rect 17 51 105 131
rect 139 17 216 97
rect 250 51 304 165
rect 338 131 499 165
rect 338 51 388 131
rect 422 17 499 97
rect 533 51 583 165
rect 617 131 782 165
rect 617 51 671 131
rect 705 17 782 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 17 199 115 340 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 920 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 25 -17 59 17 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s 37 17 59 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 37 21 884 157 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 134 157 884 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 958 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 816 51 903 165 6 X
port 6 nsew signal output
rlabel locali s 831 165 903 299 6 X
port 6 nsew signal output
rlabel locali s 816 299 903 493 6 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 920 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2932682
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2925158
<< end >>
