magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 189 21 979 157
rect 30 -17 64 17
<< scnmos >>
rect 268 47 298 131
rect 354 47 384 131
rect 440 47 470 131
rect 526 47 556 131
rect 612 47 642 131
rect 698 47 728 131
rect 784 47 814 131
rect 870 47 900 131
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 248 297 278 497
rect 332 297 362 497
rect 416 297 446 497
rect 500 297 530 497
rect 584 297 614 497
rect 668 297 698 497
rect 752 297 782 497
rect 836 297 866 497
rect 920 297 950 497
rect 1004 297 1034 497
<< ndiff >>
rect 215 95 268 131
rect 215 61 223 95
rect 257 61 268 95
rect 215 47 268 61
rect 298 106 354 131
rect 298 72 309 106
rect 343 72 354 106
rect 298 47 354 72
rect 384 95 440 131
rect 384 61 395 95
rect 429 61 440 95
rect 384 47 440 61
rect 470 106 526 131
rect 470 72 481 106
rect 515 72 526 106
rect 470 47 526 72
rect 556 95 612 131
rect 556 61 567 95
rect 601 61 612 95
rect 556 47 612 61
rect 642 106 698 131
rect 642 72 653 106
rect 687 72 698 106
rect 642 47 698 72
rect 728 95 784 131
rect 728 61 739 95
rect 773 61 784 95
rect 728 47 784 61
rect 814 106 870 131
rect 814 72 825 106
rect 859 72 870 106
rect 814 47 870 72
rect 900 95 953 131
rect 900 61 911 95
rect 945 61 953 95
rect 900 47 953 61
<< pdiff >>
rect 27 478 79 497
rect 27 444 35 478
rect 69 444 79 478
rect 27 410 79 444
rect 27 376 35 410
rect 69 376 79 410
rect 27 297 79 376
rect 109 471 163 497
rect 109 437 119 471
rect 153 437 163 471
rect 109 403 163 437
rect 109 369 119 403
rect 153 369 163 403
rect 109 297 163 369
rect 193 478 248 497
rect 193 444 204 478
rect 238 444 248 478
rect 193 410 248 444
rect 193 376 204 410
rect 238 376 248 410
rect 193 297 248 376
rect 278 471 332 497
rect 278 437 288 471
rect 322 437 332 471
rect 278 383 332 437
rect 278 349 288 383
rect 322 349 332 383
rect 278 297 332 349
rect 362 478 416 497
rect 362 444 372 478
rect 406 444 416 478
rect 362 410 416 444
rect 362 376 372 410
rect 406 376 416 410
rect 362 297 416 376
rect 446 471 500 497
rect 446 437 456 471
rect 490 437 500 471
rect 446 383 500 437
rect 446 349 456 383
rect 490 349 500 383
rect 446 297 500 349
rect 530 478 584 497
rect 530 444 540 478
rect 574 444 584 478
rect 530 410 584 444
rect 530 376 540 410
rect 574 376 584 410
rect 530 297 584 376
rect 614 471 668 497
rect 614 437 624 471
rect 658 437 668 471
rect 614 383 668 437
rect 614 349 624 383
rect 658 349 668 383
rect 614 297 668 349
rect 698 478 752 497
rect 698 444 708 478
rect 742 444 752 478
rect 698 410 752 444
rect 698 376 708 410
rect 742 376 752 410
rect 698 297 752 376
rect 782 471 836 497
rect 782 437 792 471
rect 826 437 836 471
rect 782 383 836 437
rect 782 349 792 383
rect 826 349 836 383
rect 782 297 836 349
rect 866 478 920 497
rect 866 444 876 478
rect 910 444 920 478
rect 866 410 920 444
rect 866 376 876 410
rect 910 376 920 410
rect 866 297 920 376
rect 950 471 1004 497
rect 950 437 960 471
rect 994 437 1004 471
rect 950 383 1004 437
rect 950 349 960 383
rect 994 349 1004 383
rect 950 297 1004 349
rect 1034 478 1086 497
rect 1034 444 1044 478
rect 1078 444 1086 478
rect 1034 410 1086 444
rect 1034 376 1044 410
rect 1078 376 1086 410
rect 1034 297 1086 376
<< ndiffc >>
rect 223 61 257 95
rect 309 72 343 106
rect 395 61 429 95
rect 481 72 515 106
rect 567 61 601 95
rect 653 72 687 106
rect 739 61 773 95
rect 825 72 859 106
rect 911 61 945 95
<< pdiffc >>
rect 35 444 69 478
rect 35 376 69 410
rect 119 437 153 471
rect 119 369 153 403
rect 204 444 238 478
rect 204 376 238 410
rect 288 437 322 471
rect 288 349 322 383
rect 372 444 406 478
rect 372 376 406 410
rect 456 437 490 471
rect 456 349 490 383
rect 540 444 574 478
rect 540 376 574 410
rect 624 437 658 471
rect 624 349 658 383
rect 708 444 742 478
rect 708 376 742 410
rect 792 437 826 471
rect 792 349 826 383
rect 876 444 910 478
rect 876 376 910 410
rect 960 437 994 471
rect 960 349 994 383
rect 1044 444 1078 478
rect 1044 376 1078 410
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 248 497 278 523
rect 332 497 362 523
rect 416 497 446 523
rect 500 497 530 523
rect 584 497 614 523
rect 668 497 698 523
rect 752 497 782 523
rect 836 497 866 523
rect 920 497 950 523
rect 1004 497 1034 523
rect 79 277 109 297
rect 163 277 193 297
rect 248 277 278 297
rect 332 277 362 297
rect 416 277 446 297
rect 500 277 530 297
rect 584 277 614 297
rect 668 277 698 297
rect 752 277 782 297
rect 836 277 866 297
rect 920 277 950 297
rect 1004 277 1034 297
rect 79 249 1034 277
rect 79 215 107 249
rect 141 215 175 249
rect 209 215 243 249
rect 277 215 311 249
rect 345 215 379 249
rect 413 215 447 249
rect 481 215 515 249
rect 549 215 583 249
rect 617 215 651 249
rect 685 215 719 249
rect 753 215 787 249
rect 821 215 855 249
rect 889 215 923 249
rect 957 215 1034 249
rect 79 162 1034 215
rect 268 131 298 162
rect 354 131 384 162
rect 440 131 470 162
rect 526 131 556 162
rect 612 131 642 162
rect 698 131 728 162
rect 784 131 814 162
rect 870 131 900 162
rect 268 21 298 47
rect 354 21 384 47
rect 440 21 470 47
rect 526 21 556 47
rect 612 21 642 47
rect 698 21 728 47
rect 784 21 814 47
rect 870 21 900 47
<< polycont >>
rect 107 215 141 249
rect 175 215 209 249
rect 243 215 277 249
rect 311 215 345 249
rect 379 215 413 249
rect 447 215 481 249
rect 515 215 549 249
rect 583 215 617 249
rect 651 215 685 249
rect 719 215 753 249
rect 787 215 821 249
rect 855 215 889 249
rect 923 215 957 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 27 478 79 527
rect 27 444 35 478
rect 69 444 79 478
rect 27 410 79 444
rect 27 376 35 410
rect 69 376 79 410
rect 27 360 79 376
rect 113 471 161 487
rect 113 437 119 471
rect 153 437 161 471
rect 113 403 161 437
rect 113 369 119 403
rect 153 369 161 403
rect 113 326 161 369
rect 195 478 247 527
rect 195 444 204 478
rect 238 444 247 478
rect 195 410 247 444
rect 195 376 204 410
rect 238 376 247 410
rect 195 360 247 376
rect 281 471 329 487
rect 281 437 288 471
rect 322 437 329 471
rect 281 383 329 437
rect 281 349 288 383
rect 322 349 329 383
rect 363 478 415 527
rect 363 444 372 478
rect 406 444 415 478
rect 363 410 415 444
rect 363 376 372 410
rect 406 376 415 410
rect 363 360 415 376
rect 449 471 499 487
rect 449 437 456 471
rect 490 437 499 471
rect 449 383 499 437
rect 281 326 329 349
rect 449 349 456 383
rect 490 349 499 383
rect 533 478 582 527
rect 533 444 540 478
rect 574 444 582 478
rect 533 410 582 444
rect 533 376 540 410
rect 574 376 582 410
rect 533 360 582 376
rect 616 471 665 487
rect 616 437 624 471
rect 658 437 665 471
rect 616 383 665 437
rect 449 326 499 349
rect 616 349 624 383
rect 658 349 665 383
rect 699 478 750 527
rect 699 444 708 478
rect 742 444 750 478
rect 699 410 750 444
rect 699 376 708 410
rect 742 376 750 410
rect 699 360 750 376
rect 784 471 835 487
rect 784 437 792 471
rect 826 437 835 471
rect 784 383 835 437
rect 616 326 665 349
rect 784 349 792 383
rect 826 349 835 383
rect 869 478 919 527
rect 869 444 876 478
rect 910 444 919 478
rect 869 410 919 444
rect 869 376 876 410
rect 910 376 919 410
rect 869 360 919 376
rect 953 471 1001 487
rect 953 437 960 471
rect 994 437 1001 471
rect 953 383 1001 437
rect 784 326 835 349
rect 953 349 960 383
rect 994 349 1001 383
rect 1035 478 1086 527
rect 1035 444 1044 478
rect 1078 444 1086 478
rect 1035 410 1086 444
rect 1035 376 1044 410
rect 1078 376 1086 410
rect 1035 360 1086 376
rect 953 326 1001 349
rect 23 292 1088 326
rect 23 173 57 292
rect 91 249 973 258
rect 91 215 107 249
rect 141 215 175 249
rect 209 215 243 249
rect 277 215 311 249
rect 345 215 379 249
rect 413 215 447 249
rect 481 215 515 249
rect 549 215 583 249
rect 617 215 651 249
rect 685 215 719 249
rect 753 215 787 249
rect 821 215 855 249
rect 889 215 923 249
rect 957 215 973 249
rect 91 207 973 215
rect 1034 173 1088 292
rect 23 139 1088 173
rect 307 106 345 139
rect 207 95 273 105
rect 207 61 223 95
rect 257 61 273 95
rect 207 17 273 61
rect 307 72 309 106
rect 343 72 345 106
rect 479 106 517 139
rect 307 56 345 72
rect 379 95 445 105
rect 379 61 395 95
rect 429 61 445 95
rect 379 17 445 61
rect 479 72 481 106
rect 515 72 517 106
rect 651 106 689 139
rect 479 56 517 72
rect 551 95 617 105
rect 551 61 567 95
rect 601 61 617 95
rect 551 17 617 61
rect 651 72 653 106
rect 687 72 689 106
rect 823 106 861 139
rect 651 56 689 72
rect 723 95 789 105
rect 723 61 739 95
rect 773 61 789 95
rect 723 17 789 61
rect 823 72 825 106
rect 859 72 861 106
rect 823 56 861 72
rect 895 95 961 105
rect 895 61 911 95
rect 945 61 961 95
rect 895 17 961 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 1042 289 1076 323 0 FreeSans 400 0 0 0 Y
port 6 nsew signal output
flabel locali s 1042 221 1076 255 0 FreeSans 400 0 0 0 Y
port 6 nsew signal output
flabel locali s 1042 153 1076 187 0 FreeSans 400 0 0 0 Y
port 6 nsew signal output
flabel locali s 490 221 524 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 398 221 432 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 858 221 892 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 766 221 800 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 674 221 708 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 clkinv_8
rlabel metal1 s 0 -48 1196 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1196 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_END 3359238
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3350048
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 29.900 0.000 
<< end >>
