magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< pwell >>
rect 10 76 526 1138
<< nmoslvt >>
rect 204 102 240 1112
rect 296 102 332 1112
<< ndiff >>
rect 148 1100 204 1112
rect 148 1066 159 1100
rect 193 1066 204 1100
rect 148 1032 204 1066
rect 148 998 159 1032
rect 193 998 204 1032
rect 148 964 204 998
rect 148 930 159 964
rect 193 930 204 964
rect 148 896 204 930
rect 148 862 159 896
rect 193 862 204 896
rect 148 828 204 862
rect 148 794 159 828
rect 193 794 204 828
rect 148 760 204 794
rect 148 726 159 760
rect 193 726 204 760
rect 148 692 204 726
rect 148 658 159 692
rect 193 658 204 692
rect 148 624 204 658
rect 148 590 159 624
rect 193 590 204 624
rect 148 556 204 590
rect 148 522 159 556
rect 193 522 204 556
rect 148 488 204 522
rect 148 454 159 488
rect 193 454 204 488
rect 148 420 204 454
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 240 1100 296 1112
rect 240 1066 251 1100
rect 285 1066 296 1100
rect 240 1032 296 1066
rect 240 998 251 1032
rect 285 998 296 1032
rect 240 964 296 998
rect 240 930 251 964
rect 285 930 296 964
rect 240 896 296 930
rect 240 862 251 896
rect 285 862 296 896
rect 240 828 296 862
rect 240 794 251 828
rect 285 794 296 828
rect 240 760 296 794
rect 240 726 251 760
rect 285 726 296 760
rect 240 692 296 726
rect 240 658 251 692
rect 285 658 296 692
rect 240 624 296 658
rect 240 590 251 624
rect 285 590 296 624
rect 240 556 296 590
rect 240 522 251 556
rect 285 522 296 556
rect 240 488 296 522
rect 240 454 251 488
rect 285 454 296 488
rect 240 420 296 454
rect 240 386 251 420
rect 285 386 296 420
rect 240 352 296 386
rect 240 318 251 352
rect 285 318 296 352
rect 240 284 296 318
rect 240 250 251 284
rect 285 250 296 284
rect 240 216 296 250
rect 240 182 251 216
rect 285 182 296 216
rect 240 148 296 182
rect 240 114 251 148
rect 285 114 296 148
rect 240 102 296 114
rect 332 1100 388 1112
rect 332 1066 343 1100
rect 377 1066 388 1100
rect 332 1032 388 1066
rect 332 998 343 1032
rect 377 998 388 1032
rect 332 964 388 998
rect 332 930 343 964
rect 377 930 388 964
rect 332 896 388 930
rect 332 862 343 896
rect 377 862 388 896
rect 332 828 388 862
rect 332 794 343 828
rect 377 794 388 828
rect 332 760 388 794
rect 332 726 343 760
rect 377 726 388 760
rect 332 692 388 726
rect 332 658 343 692
rect 377 658 388 692
rect 332 624 388 658
rect 332 590 343 624
rect 377 590 388 624
rect 332 556 388 590
rect 332 522 343 556
rect 377 522 388 556
rect 332 488 388 522
rect 332 454 343 488
rect 377 454 388 488
rect 332 420 388 454
rect 332 386 343 420
rect 377 386 388 420
rect 332 352 388 386
rect 332 318 343 352
rect 377 318 388 352
rect 332 284 388 318
rect 332 250 343 284
rect 377 250 388 284
rect 332 216 388 250
rect 332 182 343 216
rect 377 182 388 216
rect 332 148 388 182
rect 332 114 343 148
rect 377 114 388 148
rect 332 102 388 114
<< ndiffc >>
rect 159 1066 193 1100
rect 159 998 193 1032
rect 159 930 193 964
rect 159 862 193 896
rect 159 794 193 828
rect 159 726 193 760
rect 159 658 193 692
rect 159 590 193 624
rect 159 522 193 556
rect 159 454 193 488
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 251 1066 285 1100
rect 251 998 285 1032
rect 251 930 285 964
rect 251 862 285 896
rect 251 794 285 828
rect 251 726 285 760
rect 251 658 285 692
rect 251 590 285 624
rect 251 522 285 556
rect 251 454 285 488
rect 251 386 285 420
rect 251 318 285 352
rect 251 250 285 284
rect 251 182 285 216
rect 251 114 285 148
rect 343 1066 377 1100
rect 343 998 377 1032
rect 343 930 377 964
rect 343 862 377 896
rect 343 794 377 828
rect 343 726 377 760
rect 343 658 377 692
rect 343 590 377 624
rect 343 522 377 556
rect 343 454 377 488
rect 343 386 377 420
rect 343 318 377 352
rect 343 250 377 284
rect 343 182 377 216
rect 343 114 377 148
<< psubdiff >>
rect 36 1066 94 1112
rect 36 1032 48 1066
rect 82 1032 94 1066
rect 36 998 94 1032
rect 36 964 48 998
rect 82 964 94 998
rect 36 930 94 964
rect 36 896 48 930
rect 82 896 94 930
rect 36 862 94 896
rect 36 828 48 862
rect 82 828 94 862
rect 36 794 94 828
rect 36 760 48 794
rect 82 760 94 794
rect 36 726 94 760
rect 36 692 48 726
rect 82 692 94 726
rect 36 658 94 692
rect 36 624 48 658
rect 82 624 94 658
rect 36 590 94 624
rect 36 556 48 590
rect 82 556 94 590
rect 36 522 94 556
rect 36 488 48 522
rect 82 488 94 522
rect 36 454 94 488
rect 36 420 48 454
rect 82 420 94 454
rect 36 386 94 420
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 442 1066 500 1112
rect 442 1032 454 1066
rect 488 1032 500 1066
rect 442 998 500 1032
rect 442 964 454 998
rect 488 964 500 998
rect 442 930 500 964
rect 442 896 454 930
rect 488 896 500 930
rect 442 862 500 896
rect 442 828 454 862
rect 488 828 500 862
rect 442 794 500 828
rect 442 760 454 794
rect 488 760 500 794
rect 442 726 500 760
rect 442 692 454 726
rect 488 692 500 726
rect 442 658 500 692
rect 442 624 454 658
rect 488 624 500 658
rect 442 590 500 624
rect 442 556 454 590
rect 488 556 500 590
rect 442 522 500 556
rect 442 488 454 522
rect 488 488 500 522
rect 442 454 500 488
rect 442 420 454 454
rect 488 420 500 454
rect 442 386 500 420
rect 442 352 454 386
rect 488 352 500 386
rect 442 318 500 352
rect 442 284 454 318
rect 488 284 500 318
rect 442 250 500 284
rect 442 216 454 250
rect 488 216 500 250
rect 442 182 500 216
rect 442 148 454 182
rect 488 148 500 182
rect 442 102 500 148
<< psubdiffcont >>
rect 48 1032 82 1066
rect 48 964 82 998
rect 48 896 82 930
rect 48 828 82 862
rect 48 760 82 794
rect 48 692 82 726
rect 48 624 82 658
rect 48 556 82 590
rect 48 488 82 522
rect 48 420 82 454
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 454 1032 488 1066
rect 454 964 488 998
rect 454 896 488 930
rect 454 828 488 862
rect 454 760 488 794
rect 454 692 488 726
rect 454 624 488 658
rect 454 556 488 590
rect 454 488 488 522
rect 454 420 488 454
rect 454 352 488 386
rect 454 284 488 318
rect 454 216 488 250
rect 454 148 488 182
<< poly >>
rect 167 1184 369 1204
rect 167 1150 183 1184
rect 217 1150 251 1184
rect 285 1150 319 1184
rect 353 1150 369 1184
rect 167 1134 369 1150
rect 204 1112 240 1134
rect 296 1112 332 1134
rect 204 80 240 102
rect 296 80 332 102
rect 167 64 369 80
rect 167 30 183 64
rect 217 30 251 64
rect 285 30 319 64
rect 353 30 369 64
rect 167 10 369 30
<< polycont >>
rect 183 1150 217 1184
rect 251 1150 285 1184
rect 319 1150 353 1184
rect 183 30 217 64
rect 251 30 285 64
rect 319 30 353 64
<< locali >>
rect 167 1150 179 1184
rect 217 1150 251 1184
rect 285 1150 319 1184
rect 357 1150 369 1184
rect 159 1100 193 1116
rect 48 1020 82 1032
rect 48 948 82 964
rect 48 876 82 896
rect 48 804 82 828
rect 48 732 82 760
rect 48 660 82 692
rect 48 590 82 624
rect 48 522 82 554
rect 48 454 82 482
rect 48 386 82 410
rect 48 318 82 338
rect 48 250 82 266
rect 48 182 82 194
rect 159 1032 193 1058
rect 159 964 193 986
rect 159 896 193 914
rect 159 828 193 842
rect 159 760 193 770
rect 159 692 193 698
rect 159 624 193 626
rect 159 588 193 590
rect 159 516 193 522
rect 159 444 193 454
rect 159 372 193 386
rect 159 300 193 318
rect 159 228 193 250
rect 159 156 193 182
rect 159 98 193 114
rect 251 1100 285 1116
rect 251 1032 285 1058
rect 251 964 285 986
rect 251 896 285 914
rect 251 828 285 842
rect 251 760 285 770
rect 251 692 285 698
rect 251 624 285 626
rect 251 588 285 590
rect 251 516 285 522
rect 251 444 285 454
rect 251 372 285 386
rect 251 300 285 318
rect 251 228 285 250
rect 251 156 285 182
rect 251 98 285 114
rect 343 1100 377 1116
rect 343 1032 377 1058
rect 343 964 377 986
rect 343 896 377 914
rect 343 828 377 842
rect 343 760 377 770
rect 343 692 377 698
rect 343 624 377 626
rect 343 588 377 590
rect 343 516 377 522
rect 343 444 377 454
rect 343 372 377 386
rect 343 300 377 318
rect 343 228 377 250
rect 343 156 377 182
rect 454 1020 488 1032
rect 454 948 488 964
rect 454 876 488 896
rect 454 804 488 828
rect 454 732 488 760
rect 454 660 488 692
rect 454 590 488 624
rect 454 522 488 554
rect 454 454 488 482
rect 454 386 488 410
rect 454 318 488 338
rect 454 250 488 266
rect 454 182 488 194
rect 343 98 377 114
rect 167 30 179 64
rect 217 30 251 64
rect 285 30 319 64
rect 357 30 369 64
<< viali >>
rect 179 1150 183 1184
rect 183 1150 213 1184
rect 251 1150 285 1184
rect 323 1150 353 1184
rect 353 1150 357 1184
rect 48 1066 82 1092
rect 48 1058 82 1066
rect 48 998 82 1020
rect 48 986 82 998
rect 48 930 82 948
rect 48 914 82 930
rect 48 862 82 876
rect 48 842 82 862
rect 48 794 82 804
rect 48 770 82 794
rect 48 726 82 732
rect 48 698 82 726
rect 48 658 82 660
rect 48 626 82 658
rect 48 556 82 588
rect 48 554 82 556
rect 48 488 82 516
rect 48 482 82 488
rect 48 420 82 444
rect 48 410 82 420
rect 48 352 82 372
rect 48 338 82 352
rect 48 284 82 300
rect 48 266 82 284
rect 48 216 82 228
rect 48 194 82 216
rect 48 148 82 156
rect 48 122 82 148
rect 159 1066 193 1092
rect 159 1058 193 1066
rect 159 998 193 1020
rect 159 986 193 998
rect 159 930 193 948
rect 159 914 193 930
rect 159 862 193 876
rect 159 842 193 862
rect 159 794 193 804
rect 159 770 193 794
rect 159 726 193 732
rect 159 698 193 726
rect 159 658 193 660
rect 159 626 193 658
rect 159 556 193 588
rect 159 554 193 556
rect 159 488 193 516
rect 159 482 193 488
rect 159 420 193 444
rect 159 410 193 420
rect 159 352 193 372
rect 159 338 193 352
rect 159 284 193 300
rect 159 266 193 284
rect 159 216 193 228
rect 159 194 193 216
rect 159 148 193 156
rect 159 122 193 148
rect 251 1066 285 1092
rect 251 1058 285 1066
rect 251 998 285 1020
rect 251 986 285 998
rect 251 930 285 948
rect 251 914 285 930
rect 251 862 285 876
rect 251 842 285 862
rect 251 794 285 804
rect 251 770 285 794
rect 251 726 285 732
rect 251 698 285 726
rect 251 658 285 660
rect 251 626 285 658
rect 251 556 285 588
rect 251 554 285 556
rect 251 488 285 516
rect 251 482 285 488
rect 251 420 285 444
rect 251 410 285 420
rect 251 352 285 372
rect 251 338 285 352
rect 251 284 285 300
rect 251 266 285 284
rect 251 216 285 228
rect 251 194 285 216
rect 251 148 285 156
rect 251 122 285 148
rect 343 1066 377 1092
rect 343 1058 377 1066
rect 343 998 377 1020
rect 343 986 377 998
rect 343 930 377 948
rect 343 914 377 930
rect 343 862 377 876
rect 343 842 377 862
rect 343 794 377 804
rect 343 770 377 794
rect 343 726 377 732
rect 343 698 377 726
rect 343 658 377 660
rect 343 626 377 658
rect 343 556 377 588
rect 343 554 377 556
rect 343 488 377 516
rect 343 482 377 488
rect 343 420 377 444
rect 343 410 377 420
rect 343 352 377 372
rect 343 338 377 352
rect 343 284 377 300
rect 343 266 377 284
rect 343 216 377 228
rect 343 194 377 216
rect 343 148 377 156
rect 343 122 377 148
rect 454 1066 488 1092
rect 454 1058 488 1066
rect 454 998 488 1020
rect 454 986 488 998
rect 454 930 488 948
rect 454 914 488 930
rect 454 862 488 876
rect 454 842 488 862
rect 454 794 488 804
rect 454 770 488 794
rect 454 726 488 732
rect 454 698 488 726
rect 454 658 488 660
rect 454 626 488 658
rect 454 556 488 588
rect 454 554 488 556
rect 454 488 488 516
rect 454 482 488 488
rect 454 420 488 444
rect 454 410 488 420
rect 454 352 488 372
rect 454 338 488 352
rect 454 284 488 300
rect 454 266 488 284
rect 454 216 488 228
rect 454 194 488 216
rect 454 148 488 156
rect 454 122 488 148
rect 179 30 183 64
rect 183 30 213 64
rect 251 30 285 64
rect 323 30 353 64
rect 353 30 357 64
<< metal1 >>
rect 167 1184 369 1204
rect 167 1150 179 1184
rect 213 1150 251 1184
rect 285 1150 323 1184
rect 357 1150 369 1184
rect 167 1138 369 1150
rect 36 1092 94 1104
rect 36 1058 48 1092
rect 82 1058 94 1092
rect 36 1020 94 1058
rect 36 986 48 1020
rect 82 986 94 1020
rect 36 948 94 986
rect 36 914 48 948
rect 82 914 94 948
rect 36 876 94 914
rect 36 842 48 876
rect 82 842 94 876
rect 36 804 94 842
rect 36 770 48 804
rect 82 770 94 804
rect 36 732 94 770
rect 36 698 48 732
rect 82 698 94 732
rect 36 660 94 698
rect 36 626 48 660
rect 82 626 94 660
rect 36 588 94 626
rect 36 554 48 588
rect 82 554 94 588
rect 36 516 94 554
rect 36 482 48 516
rect 82 482 94 516
rect 36 444 94 482
rect 36 410 48 444
rect 82 410 94 444
rect 36 372 94 410
rect 36 338 48 372
rect 82 338 94 372
rect 36 300 94 338
rect 36 266 48 300
rect 82 266 94 300
rect 36 228 94 266
rect 36 194 48 228
rect 82 194 94 228
rect 36 156 94 194
rect 36 122 48 156
rect 82 122 94 156
rect 36 110 94 122
rect 150 1092 202 1104
rect 150 1058 159 1092
rect 193 1058 202 1092
rect 150 1020 202 1058
rect 150 986 159 1020
rect 193 986 202 1020
rect 150 948 202 986
rect 150 914 159 948
rect 193 914 202 948
rect 150 876 202 914
rect 150 842 159 876
rect 193 842 202 876
rect 150 804 202 842
rect 150 770 159 804
rect 193 770 202 804
rect 150 732 202 770
rect 150 698 159 732
rect 193 698 202 732
rect 150 660 202 698
rect 150 626 159 660
rect 193 626 202 660
rect 150 588 202 626
rect 150 554 159 588
rect 193 554 202 588
rect 150 552 202 554
rect 150 488 159 500
rect 193 488 202 500
rect 150 424 159 436
rect 193 424 202 436
rect 150 360 159 372
rect 193 360 202 372
rect 150 300 202 308
rect 150 296 159 300
rect 193 296 202 300
rect 150 232 202 244
rect 150 168 202 180
rect 150 110 202 116
rect 242 1098 294 1104
rect 242 1034 294 1046
rect 242 970 294 982
rect 242 914 251 918
rect 285 914 294 918
rect 242 906 294 914
rect 242 842 251 854
rect 285 842 294 854
rect 242 778 251 790
rect 285 778 294 790
rect 242 714 251 726
rect 285 714 294 726
rect 242 660 294 662
rect 242 626 251 660
rect 285 626 294 660
rect 242 588 294 626
rect 242 554 251 588
rect 285 554 294 588
rect 242 516 294 554
rect 242 482 251 516
rect 285 482 294 516
rect 242 444 294 482
rect 242 410 251 444
rect 285 410 294 444
rect 242 372 294 410
rect 242 338 251 372
rect 285 338 294 372
rect 242 300 294 338
rect 242 266 251 300
rect 285 266 294 300
rect 242 228 294 266
rect 242 194 251 228
rect 285 194 294 228
rect 242 156 294 194
rect 242 122 251 156
rect 285 122 294 156
rect 242 110 294 122
rect 334 1092 386 1104
rect 334 1058 343 1092
rect 377 1058 386 1092
rect 334 1020 386 1058
rect 334 986 343 1020
rect 377 986 386 1020
rect 334 948 386 986
rect 334 914 343 948
rect 377 914 386 948
rect 334 876 386 914
rect 334 842 343 876
rect 377 842 386 876
rect 334 804 386 842
rect 334 770 343 804
rect 377 770 386 804
rect 334 732 386 770
rect 334 698 343 732
rect 377 698 386 732
rect 334 660 386 698
rect 334 626 343 660
rect 377 626 386 660
rect 334 588 386 626
rect 334 554 343 588
rect 377 554 386 588
rect 334 552 386 554
rect 334 488 343 500
rect 377 488 386 500
rect 334 424 343 436
rect 377 424 386 436
rect 334 360 343 372
rect 377 360 386 372
rect 334 300 386 308
rect 334 296 343 300
rect 377 296 386 300
rect 334 232 386 244
rect 334 168 386 180
rect 334 110 386 116
rect 442 1092 500 1104
rect 442 1058 454 1092
rect 488 1058 500 1092
rect 442 1020 500 1058
rect 442 986 454 1020
rect 488 986 500 1020
rect 442 948 500 986
rect 442 914 454 948
rect 488 914 500 948
rect 442 876 500 914
rect 442 842 454 876
rect 488 842 500 876
rect 442 804 500 842
rect 442 770 454 804
rect 488 770 500 804
rect 442 732 500 770
rect 442 698 454 732
rect 488 698 500 732
rect 442 660 500 698
rect 442 626 454 660
rect 488 626 500 660
rect 442 588 500 626
rect 442 554 454 588
rect 488 554 500 588
rect 442 516 500 554
rect 442 482 454 516
rect 488 482 500 516
rect 442 444 500 482
rect 442 410 454 444
rect 488 410 500 444
rect 442 372 500 410
rect 442 338 454 372
rect 488 338 500 372
rect 442 300 500 338
rect 442 266 454 300
rect 488 266 500 300
rect 442 228 500 266
rect 442 194 454 228
rect 488 194 500 228
rect 442 156 500 194
rect 442 122 454 156
rect 488 122 500 156
rect 442 110 500 122
rect 167 64 369 76
rect 167 30 179 64
rect 213 30 251 64
rect 285 30 323 64
rect 357 30 369 64
rect 167 10 369 30
<< via1 >>
rect 150 516 202 552
rect 150 500 159 516
rect 159 500 193 516
rect 193 500 202 516
rect 150 482 159 488
rect 159 482 193 488
rect 193 482 202 488
rect 150 444 202 482
rect 150 436 159 444
rect 159 436 193 444
rect 193 436 202 444
rect 150 410 159 424
rect 159 410 193 424
rect 193 410 202 424
rect 150 372 202 410
rect 150 338 159 360
rect 159 338 193 360
rect 193 338 202 360
rect 150 308 202 338
rect 150 266 159 296
rect 159 266 193 296
rect 193 266 202 296
rect 150 244 202 266
rect 150 228 202 232
rect 150 194 159 228
rect 159 194 193 228
rect 193 194 202 228
rect 150 180 202 194
rect 150 156 202 168
rect 150 122 159 156
rect 159 122 193 156
rect 193 122 202 156
rect 150 116 202 122
rect 242 1092 294 1098
rect 242 1058 251 1092
rect 251 1058 285 1092
rect 285 1058 294 1092
rect 242 1046 294 1058
rect 242 1020 294 1034
rect 242 986 251 1020
rect 251 986 285 1020
rect 285 986 294 1020
rect 242 982 294 986
rect 242 948 294 970
rect 242 918 251 948
rect 251 918 285 948
rect 285 918 294 948
rect 242 876 294 906
rect 242 854 251 876
rect 251 854 285 876
rect 285 854 294 876
rect 242 804 294 842
rect 242 790 251 804
rect 251 790 285 804
rect 285 790 294 804
rect 242 770 251 778
rect 251 770 285 778
rect 285 770 294 778
rect 242 732 294 770
rect 242 726 251 732
rect 251 726 285 732
rect 285 726 294 732
rect 242 698 251 714
rect 251 698 285 714
rect 285 698 294 714
rect 242 662 294 698
rect 334 516 386 552
rect 334 500 343 516
rect 343 500 377 516
rect 377 500 386 516
rect 334 482 343 488
rect 343 482 377 488
rect 377 482 386 488
rect 334 444 386 482
rect 334 436 343 444
rect 343 436 377 444
rect 377 436 386 444
rect 334 410 343 424
rect 343 410 377 424
rect 377 410 386 424
rect 334 372 386 410
rect 334 338 343 360
rect 343 338 377 360
rect 377 338 386 360
rect 334 308 386 338
rect 334 266 343 296
rect 343 266 377 296
rect 377 266 386 296
rect 334 244 386 266
rect 334 228 386 232
rect 334 194 343 228
rect 343 194 377 228
rect 377 194 386 228
rect 334 180 386 194
rect 334 156 386 168
rect 334 122 343 156
rect 343 122 377 156
rect 377 122 386 156
rect 334 116 386 122
<< metal2 >>
rect 10 1098 526 1104
rect 10 1046 242 1098
rect 294 1046 526 1098
rect 10 1034 526 1046
rect 10 982 242 1034
rect 294 982 526 1034
rect 10 970 526 982
rect 10 918 242 970
rect 294 918 526 970
rect 10 906 526 918
rect 10 854 242 906
rect 294 854 526 906
rect 10 842 526 854
rect 10 790 242 842
rect 294 790 526 842
rect 10 778 526 790
rect 10 726 242 778
rect 294 726 526 778
rect 10 714 526 726
rect 10 662 242 714
rect 294 662 526 714
rect 10 632 526 662
rect 10 552 526 582
rect 10 500 150 552
rect 202 500 334 552
rect 386 500 526 552
rect 10 488 526 500
rect 10 436 150 488
rect 202 436 334 488
rect 386 436 526 488
rect 10 424 526 436
rect 10 372 150 424
rect 202 372 334 424
rect 386 372 526 424
rect 10 360 526 372
rect 10 308 150 360
rect 202 308 334 360
rect 386 308 526 360
rect 10 296 526 308
rect 10 244 150 296
rect 202 244 334 296
rect 386 244 526 296
rect 10 232 526 244
rect 10 180 150 232
rect 202 180 334 232
rect 386 180 526 232
rect 10 168 526 180
rect 10 116 150 168
rect 202 116 334 168
rect 386 116 526 168
rect 10 110 526 116
<< labels >>
flabel metal2 s 10 632 30 1104 7 FreeSans 300 180 0 0 DRAIN
port 2 nsew
flabel metal2 s 10 110 30 582 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal1 s 167 1138 369 1204 0 FreeSans 300 0 0 0 GATE
port 4 nsew
flabel metal1 s 167 10 369 76 0 FreeSans 300 0 0 0 GATE
port 4 nsew
flabel metal1 s 442 110 500 126 3 FreeSans 300 90 0 0 SUBSTRATE
port 5 nsew
flabel metal1 s 36 110 94 126 3 FreeSans 300 90 0 0 SUBSTRATE
port 5 nsew
<< properties >>
string GDS_END 5960942
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 5945470
<< end >>
