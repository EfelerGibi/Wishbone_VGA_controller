magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -66 377 1026 897
<< pwell >>
rect 66 43 956 283
rect -26 -43 986 43
<< mvnmos >>
rect 149 107 249 257
rect 305 107 405 257
rect 461 107 561 257
rect 617 107 717 257
rect 773 107 873 257
<< mvpmos >>
rect 149 443 249 743
rect 305 443 405 743
rect 461 443 561 743
rect 617 443 717 743
rect 773 443 873 743
<< mvndiff >>
rect 92 249 149 257
rect 92 215 104 249
rect 138 215 149 249
rect 92 149 149 215
rect 92 115 104 149
rect 138 115 149 149
rect 92 107 149 115
rect 249 249 305 257
rect 249 215 260 249
rect 294 215 305 249
rect 249 149 305 215
rect 249 115 260 149
rect 294 115 305 149
rect 249 107 305 115
rect 405 177 461 257
rect 405 143 416 177
rect 450 143 461 177
rect 405 107 461 143
rect 561 249 617 257
rect 561 215 572 249
rect 606 215 617 249
rect 561 149 617 215
rect 561 115 572 149
rect 606 115 617 149
rect 561 107 617 115
rect 717 249 773 257
rect 717 215 728 249
rect 762 215 773 249
rect 717 149 773 215
rect 717 115 728 149
rect 762 115 773 149
rect 717 107 773 115
rect 873 249 930 257
rect 873 215 884 249
rect 918 215 930 249
rect 873 149 930 215
rect 873 115 884 149
rect 918 115 930 149
rect 873 107 930 115
<< mvpdiff >>
rect 92 735 149 743
rect 92 701 104 735
rect 138 701 149 735
rect 92 652 149 701
rect 92 618 104 652
rect 138 618 149 652
rect 92 568 149 618
rect 92 534 104 568
rect 138 534 149 568
rect 92 485 149 534
rect 92 451 104 485
rect 138 451 149 485
rect 92 443 149 451
rect 249 735 305 743
rect 249 701 260 735
rect 294 701 305 735
rect 249 652 305 701
rect 249 618 260 652
rect 294 618 305 652
rect 249 568 305 618
rect 249 534 260 568
rect 294 534 305 568
rect 249 485 305 534
rect 249 451 260 485
rect 294 451 305 485
rect 249 443 305 451
rect 405 735 461 743
rect 405 701 416 735
rect 450 701 461 735
rect 405 652 461 701
rect 405 618 416 652
rect 450 618 461 652
rect 405 568 461 618
rect 405 534 416 568
rect 450 534 461 568
rect 405 485 461 534
rect 405 451 416 485
rect 450 451 461 485
rect 405 443 461 451
rect 561 735 617 743
rect 561 701 572 735
rect 606 701 617 735
rect 561 652 617 701
rect 561 618 572 652
rect 606 618 617 652
rect 561 568 617 618
rect 561 534 572 568
rect 606 534 617 568
rect 561 485 617 534
rect 561 451 572 485
rect 606 451 617 485
rect 561 443 617 451
rect 717 735 773 743
rect 717 701 728 735
rect 762 701 773 735
rect 717 655 773 701
rect 717 621 728 655
rect 762 621 773 655
rect 717 574 773 621
rect 717 540 728 574
rect 762 540 773 574
rect 717 494 773 540
rect 717 460 728 494
rect 762 460 773 494
rect 717 443 773 460
rect 873 735 930 743
rect 873 701 884 735
rect 918 701 930 735
rect 873 652 930 701
rect 873 618 884 652
rect 918 618 930 652
rect 873 568 930 618
rect 873 534 884 568
rect 918 534 930 568
rect 873 485 930 534
rect 873 451 884 485
rect 918 451 930 485
rect 873 443 930 451
<< mvndiffc >>
rect 104 215 138 249
rect 104 115 138 149
rect 260 215 294 249
rect 260 115 294 149
rect 416 143 450 177
rect 572 215 606 249
rect 572 115 606 149
rect 728 215 762 249
rect 728 115 762 149
rect 884 215 918 249
rect 884 115 918 149
<< mvpdiffc >>
rect 104 701 138 735
rect 104 618 138 652
rect 104 534 138 568
rect 104 451 138 485
rect 260 701 294 735
rect 260 618 294 652
rect 260 534 294 568
rect 260 451 294 485
rect 416 701 450 735
rect 416 618 450 652
rect 416 534 450 568
rect 416 451 450 485
rect 572 701 606 735
rect 572 618 606 652
rect 572 534 606 568
rect 572 451 606 485
rect 728 701 762 735
rect 728 621 762 655
rect 728 540 762 574
rect 728 460 762 494
rect 884 701 918 735
rect 884 618 918 652
rect 884 534 918 568
rect 884 451 918 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 960 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
<< poly >>
rect 149 743 249 769
rect 305 743 405 769
rect 461 743 561 769
rect 617 743 717 769
rect 773 743 873 769
rect 149 383 249 443
rect 305 383 405 443
rect 461 383 561 443
rect 617 383 717 443
rect 773 395 873 443
rect 149 345 724 383
rect 149 311 330 345
rect 364 311 398 345
rect 432 311 466 345
rect 500 311 534 345
rect 568 311 602 345
rect 636 311 670 345
rect 704 311 724 345
rect 149 283 724 311
rect 773 361 793 395
rect 827 361 873 395
rect 149 257 249 283
rect 305 257 405 283
rect 461 257 561 283
rect 617 257 717 283
rect 773 257 873 361
rect 149 81 249 107
rect 305 81 405 107
rect 461 81 561 107
rect 617 81 717 107
rect 773 81 873 107
<< polycont >>
rect 330 311 364 345
rect 398 311 432 345
rect 466 311 500 345
rect 534 311 568 345
rect 602 311 636 345
rect 670 311 704 345
rect 793 361 827 395
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 960 831
rect 18 735 208 751
rect 18 701 24 735
rect 58 701 96 735
rect 138 701 168 735
rect 202 701 208 735
rect 18 652 208 701
rect 18 618 104 652
rect 138 618 208 652
rect 18 568 208 618
rect 18 534 104 568
rect 138 534 208 568
rect 18 485 208 534
rect 18 451 104 485
rect 138 451 208 485
rect 18 435 208 451
rect 244 735 294 751
rect 244 701 260 735
rect 244 652 294 701
rect 244 618 260 652
rect 244 568 294 618
rect 244 534 260 568
rect 244 485 294 534
rect 244 451 260 485
rect 330 735 520 751
rect 330 701 336 735
rect 370 701 408 735
rect 450 701 480 735
rect 514 701 520 735
rect 330 652 520 701
rect 330 618 416 652
rect 450 618 520 652
rect 330 568 520 618
rect 330 534 416 568
rect 450 534 520 568
rect 330 485 520 534
rect 330 451 416 485
rect 450 451 520 485
rect 556 735 622 751
rect 556 701 572 735
rect 606 701 622 735
rect 556 652 622 701
rect 556 618 572 652
rect 606 618 622 652
rect 556 568 622 618
rect 556 534 572 568
rect 606 534 622 568
rect 556 485 622 534
rect 556 451 572 485
rect 606 451 622 485
rect 658 735 848 751
rect 658 701 664 735
rect 698 701 728 735
rect 770 701 808 735
rect 842 701 848 735
rect 658 655 848 701
rect 658 621 728 655
rect 762 621 848 655
rect 658 574 848 621
rect 658 540 728 574
rect 762 540 848 574
rect 658 494 848 540
rect 658 460 728 494
rect 762 460 848 494
rect 884 735 934 751
rect 918 701 934 735
rect 884 652 934 701
rect 918 618 934 652
rect 884 568 934 618
rect 918 534 934 568
rect 884 485 934 534
rect 244 415 294 451
rect 556 415 622 451
rect 918 451 934 485
rect 244 381 622 415
rect 777 395 843 424
rect 244 356 278 381
rect 25 310 278 356
rect 777 361 793 395
rect 827 361 843 395
rect 777 355 843 361
rect 314 311 330 345
rect 364 311 398 345
rect 432 311 466 345
rect 500 311 534 345
rect 568 311 602 345
rect 636 311 670 345
rect 704 319 720 345
rect 884 319 934 451
rect 704 311 934 319
rect 244 275 278 310
rect 686 285 934 311
rect 18 249 208 265
rect 18 215 104 249
rect 138 215 208 249
rect 18 149 208 215
rect 18 115 104 149
rect 138 115 208 149
rect 18 113 208 115
rect 18 79 24 113
rect 58 79 96 113
rect 130 79 168 113
rect 202 79 208 113
rect 244 249 606 275
rect 868 249 934 285
rect 244 215 260 249
rect 294 241 572 249
rect 244 149 294 215
rect 556 215 572 241
rect 244 115 260 149
rect 244 99 294 115
rect 330 177 520 205
rect 330 143 416 177
rect 450 143 520 177
rect 330 113 520 143
rect 18 73 208 79
rect 330 79 336 113
rect 370 79 408 113
rect 442 79 480 113
rect 514 79 520 113
rect 556 149 606 215
rect 556 115 572 149
rect 556 99 606 115
rect 642 215 728 249
rect 762 215 832 249
rect 642 149 832 215
rect 642 115 728 149
rect 762 115 832 149
rect 642 113 832 115
rect 330 73 520 79
rect 642 79 648 113
rect 682 79 720 113
rect 754 79 792 113
rect 826 79 832 113
rect 868 215 884 249
rect 918 215 934 249
rect 868 149 934 215
rect 868 115 884 149
rect 918 115 934 149
rect 868 99 934 115
rect 642 73 832 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 24 701 58 735
rect 96 701 104 735
rect 104 701 130 735
rect 168 701 202 735
rect 336 701 370 735
rect 408 701 416 735
rect 416 701 442 735
rect 480 701 514 735
rect 664 701 698 735
rect 736 701 762 735
rect 762 701 770 735
rect 808 701 842 735
rect 24 79 58 113
rect 96 79 130 113
rect 168 79 202 113
rect 336 79 370 113
rect 408 79 442 113
rect 480 79 514 113
rect 648 79 682 113
rect 720 79 754 113
rect 792 79 826 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 831 960 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 960 831
rect 0 791 960 797
rect 0 735 960 763
rect 0 701 24 735
rect 58 701 96 735
rect 130 701 168 735
rect 202 701 336 735
rect 370 701 408 735
rect 442 701 480 735
rect 514 701 664 735
rect 698 701 736 735
rect 770 701 808 735
rect 842 701 960 735
rect 0 689 960 701
rect 0 113 960 125
rect 0 79 24 113
rect 58 79 96 113
rect 130 79 168 113
rect 202 79 336 113
rect 370 79 408 113
rect 442 79 480 113
rect 514 79 648 113
rect 682 79 720 113
rect 754 79 792 113
rect 826 79 960 113
rect 0 51 960 79
rect 0 17 960 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -23 960 -17
<< labels >>
rlabel comment s 0 0 0 0 4 buf_4
flabel metal1 s 0 51 960 125 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 0 0 960 23 0 FreeSans 340 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 0 689 960 763 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 791 960 814 0 FreeSans 340 0 0 0 VPB
port 4 nsew power bidirectional
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 960 814
string GDS_END 841122
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 829916
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
