magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< metal1 >>
rect 1465 2168 1471 2220
rect 1523 2168 1529 2220
rect 1570 1130 1604 2256
rect 1646 1142 1674 2256
rect 3961 2168 3967 2220
rect 4019 2168 4025 2220
rect 1793 2016 1799 2068
rect 1851 2016 1857 2068
rect 1711 1242 1717 1294
rect 1769 1242 1775 1294
rect 4066 1130 4100 2256
rect 4142 1142 4170 2256
rect 6457 2168 6463 2220
rect 6515 2168 6521 2220
rect 4289 2016 4295 2068
rect 4347 2016 4353 2068
rect 4207 1242 4213 1294
rect 4265 1242 4271 1294
rect 6562 1130 6596 2256
rect 6638 1142 6666 2256
rect 8953 2168 8959 2220
rect 9011 2168 9017 2220
rect 6785 2016 6791 2068
rect 6843 2016 6849 2068
rect 6703 1242 6709 1294
rect 6761 1242 6767 1294
rect 9058 1130 9092 2256
rect 9134 1142 9162 2256
rect 11449 2168 11455 2220
rect 11507 2168 11513 2220
rect 9281 2016 9287 2068
rect 9339 2016 9345 2068
rect 9199 1242 9205 1294
rect 9257 1242 9263 1294
rect 11554 1130 11588 2256
rect 11630 1142 11658 2256
rect 13945 2168 13951 2220
rect 14003 2168 14009 2220
rect 11777 2016 11783 2068
rect 11835 2016 11841 2068
rect 11695 1242 11701 1294
rect 11753 1242 11759 1294
rect 14050 1130 14084 2256
rect 14126 1142 14154 2256
rect 16441 2168 16447 2220
rect 16499 2168 16505 2220
rect 14273 2016 14279 2068
rect 14331 2016 14337 2068
rect 14191 1242 14197 1294
rect 14249 1242 14255 1294
rect 16546 1130 16580 2256
rect 16622 1142 16650 2256
rect 18937 2168 18943 2220
rect 18995 2168 19001 2220
rect 16769 2016 16775 2068
rect 16827 2016 16833 2068
rect 16687 1242 16693 1294
rect 16745 1242 16751 1294
rect 19042 1130 19076 2256
rect 19118 1142 19146 2256
rect 21433 2168 21439 2220
rect 21491 2168 21497 2220
rect 19265 2016 19271 2068
rect 19323 2016 19329 2068
rect 19183 1242 19189 1294
rect 19241 1242 19247 1294
rect 21538 1130 21572 2256
rect 21614 1142 21642 2256
rect 23929 2168 23935 2220
rect 23987 2168 23993 2220
rect 21761 2016 21767 2068
rect 21819 2016 21825 2068
rect 21679 1242 21685 1294
rect 21737 1242 21743 1294
rect 24034 1130 24068 2256
rect 24110 1142 24138 2256
rect 26425 2168 26431 2220
rect 26483 2168 26489 2220
rect 24257 2016 24263 2068
rect 24315 2016 24321 2068
rect 24175 1242 24181 1294
rect 24233 1242 24239 1294
rect 26530 1130 26564 2256
rect 26606 1142 26634 2256
rect 28921 2168 28927 2220
rect 28979 2168 28985 2220
rect 26753 2016 26759 2068
rect 26811 2016 26817 2068
rect 26671 1242 26677 1294
rect 26729 1242 26735 1294
rect 29026 1130 29060 2256
rect 29102 1142 29130 2256
rect 31417 2168 31423 2220
rect 31475 2168 31481 2220
rect 29249 2016 29255 2068
rect 29307 2016 29313 2068
rect 29167 1242 29173 1294
rect 29225 1242 29231 1294
rect 31522 1130 31556 2256
rect 31598 1142 31626 2256
rect 33913 2168 33919 2220
rect 33971 2168 33977 2220
rect 31745 2016 31751 2068
rect 31803 2016 31809 2068
rect 31663 1242 31669 1294
rect 31721 1242 31727 1294
rect 34018 1130 34052 2256
rect 34094 1142 34122 2256
rect 36409 2168 36415 2220
rect 36467 2168 36473 2220
rect 34241 2016 34247 2068
rect 34299 2016 34305 2068
rect 34159 1242 34165 1294
rect 34217 1242 34223 1294
rect 36514 1130 36548 2256
rect 36590 1142 36618 2256
rect 38905 2168 38911 2220
rect 38963 2168 38969 2220
rect 36737 2016 36743 2068
rect 36795 2016 36801 2068
rect 36655 1242 36661 1294
rect 36713 1242 36719 1294
rect 39010 1130 39044 2256
rect 39086 1142 39114 2256
rect 41401 2168 41407 2220
rect 41459 2168 41465 2220
rect 39233 2016 39239 2068
rect 39291 2016 39297 2068
rect 39151 1242 39157 1294
rect 39209 1242 39215 1294
rect 41506 1130 41540 2256
rect 41582 1142 41610 2256
rect 43897 2168 43903 2220
rect 43955 2168 43961 2220
rect 41729 2016 41735 2068
rect 41787 2016 41793 2068
rect 41647 1242 41653 1294
rect 41705 1242 41711 1294
rect 44002 1130 44036 2256
rect 44078 1142 44106 2256
rect 46393 2168 46399 2220
rect 46451 2168 46457 2220
rect 44225 2016 44231 2068
rect 44283 2016 44289 2068
rect 44143 1242 44149 1294
rect 44201 1242 44207 1294
rect 46498 1130 46532 2256
rect 46574 1142 46602 2256
rect 48889 2168 48895 2220
rect 48947 2168 48953 2220
rect 46721 2016 46727 2068
rect 46779 2016 46785 2068
rect 46639 1242 46645 1294
rect 46697 1242 46703 1294
rect 48994 1130 49028 2256
rect 49070 1142 49098 2256
rect 51385 2168 51391 2220
rect 51443 2168 51449 2220
rect 49217 2016 49223 2068
rect 49275 2016 49281 2068
rect 49135 1242 49141 1294
rect 49193 1242 49199 1294
rect 51490 1130 51524 2256
rect 51566 1142 51594 2256
rect 53881 2168 53887 2220
rect 53939 2168 53945 2220
rect 51713 2016 51719 2068
rect 51771 2016 51777 2068
rect 51631 1242 51637 1294
rect 51689 1242 51695 1294
rect 53986 1130 54020 2256
rect 54062 1142 54090 2256
rect 56377 2168 56383 2220
rect 56435 2168 56441 2220
rect 54209 2016 54215 2068
rect 54267 2016 54273 2068
rect 54127 1242 54133 1294
rect 54185 1242 54191 1294
rect 56482 1130 56516 2256
rect 56558 1142 56586 2256
rect 58873 2168 58879 2220
rect 58931 2168 58937 2220
rect 56705 2016 56711 2068
rect 56763 2016 56769 2068
rect 56623 1242 56629 1294
rect 56681 1242 56687 1294
rect 58978 1130 59012 2256
rect 59054 1142 59082 2256
rect 61369 2168 61375 2220
rect 61427 2168 61433 2220
rect 59201 2016 59207 2068
rect 59259 2016 59265 2068
rect 59119 1242 59125 1294
rect 59177 1242 59183 1294
rect 61474 1130 61508 2256
rect 61550 1142 61578 2256
rect 63865 2168 63871 2220
rect 63923 2168 63929 2220
rect 61697 2016 61703 2068
rect 61755 2016 61761 2068
rect 61615 1242 61621 1294
rect 61673 1242 61679 1294
rect 63970 1130 64004 2256
rect 64046 1142 64074 2256
rect 66361 2168 66367 2220
rect 66419 2168 66425 2220
rect 64193 2016 64199 2068
rect 64251 2016 64257 2068
rect 64111 1242 64117 1294
rect 64169 1242 64175 1294
rect 66466 1130 66500 2256
rect 66542 1142 66570 2256
rect 68857 2168 68863 2220
rect 68915 2168 68921 2220
rect 66689 2016 66695 2068
rect 66747 2016 66753 2068
rect 66607 1242 66613 1294
rect 66665 1242 66671 1294
rect 68962 1130 68996 2256
rect 69038 1142 69066 2256
rect 71353 2168 71359 2220
rect 71411 2168 71417 2220
rect 69185 2016 69191 2068
rect 69243 2016 69249 2068
rect 69103 1242 69109 1294
rect 69161 1242 69167 1294
rect 71458 1130 71492 2256
rect 71534 1142 71562 2256
rect 73849 2168 73855 2220
rect 73907 2168 73913 2220
rect 71681 2016 71687 2068
rect 71739 2016 71745 2068
rect 71599 1242 71605 1294
rect 71657 1242 71663 1294
rect 73954 1130 73988 2256
rect 74030 1142 74058 2256
rect 76345 2168 76351 2220
rect 76403 2168 76409 2220
rect 74177 2016 74183 2068
rect 74235 2016 74241 2068
rect 74095 1242 74101 1294
rect 74153 1242 74159 1294
rect 76450 1130 76484 2256
rect 76526 1142 76554 2256
rect 78841 2168 78847 2220
rect 78899 2168 78905 2220
rect 76673 2016 76679 2068
rect 76731 2016 76737 2068
rect 76591 1242 76597 1294
rect 76649 1242 76655 1294
rect 78946 1130 78980 2256
rect 79022 1142 79050 2256
rect 79169 2016 79175 2068
rect 79227 2016 79233 2068
rect 79087 1242 79093 1294
rect 79145 1242 79151 1294
rect 1723 404 1729 456
rect 1781 404 1787 456
rect 4219 404 4225 456
rect 4277 404 4283 456
rect 6715 404 6721 456
rect 6773 404 6779 456
rect 9211 404 9217 456
rect 9269 404 9275 456
rect 11707 404 11713 456
rect 11765 404 11771 456
rect 14203 404 14209 456
rect 14261 404 14267 456
rect 16699 404 16705 456
rect 16757 404 16763 456
rect 19195 404 19201 456
rect 19253 404 19259 456
rect 21691 404 21697 456
rect 21749 404 21755 456
rect 24187 404 24193 456
rect 24245 404 24251 456
rect 26683 404 26689 456
rect 26741 404 26747 456
rect 29179 404 29185 456
rect 29237 404 29243 456
rect 31675 404 31681 456
rect 31733 404 31739 456
rect 34171 404 34177 456
rect 34229 404 34235 456
rect 36667 404 36673 456
rect 36725 404 36731 456
rect 39163 404 39169 456
rect 39221 404 39227 456
rect 41659 404 41665 456
rect 41717 404 41723 456
rect 44155 404 44161 456
rect 44213 404 44219 456
rect 46651 404 46657 456
rect 46709 404 46715 456
rect 49147 404 49153 456
rect 49205 404 49211 456
rect 51643 404 51649 456
rect 51701 404 51707 456
rect 54139 404 54145 456
rect 54197 404 54203 456
rect 56635 404 56641 456
rect 56693 404 56699 456
rect 59131 404 59137 456
rect 59189 404 59195 456
rect 61627 404 61633 456
rect 61685 404 61691 456
rect 64123 404 64129 456
rect 64181 404 64187 456
rect 66619 404 66625 456
rect 66677 404 66683 456
rect 69115 404 69121 456
rect 69173 404 69179 456
rect 71611 404 71617 456
rect 71669 404 71675 456
rect 74107 404 74113 456
rect 74165 404 74171 456
rect 76603 404 76609 456
rect 76661 404 76667 456
rect 79099 404 79105 456
rect 79157 404 79163 456
rect 1478 0 1524 254
rect 1723 82 1729 134
rect 1781 82 1787 134
rect 3974 0 4020 254
rect 4219 82 4225 134
rect 4277 82 4283 134
rect 6470 0 6516 254
rect 6715 82 6721 134
rect 6773 82 6779 134
rect 8966 0 9012 254
rect 9211 82 9217 134
rect 9269 82 9275 134
rect 11462 0 11508 254
rect 11707 82 11713 134
rect 11765 82 11771 134
rect 13958 0 14004 254
rect 14203 82 14209 134
rect 14261 82 14267 134
rect 16454 0 16500 254
rect 16699 82 16705 134
rect 16757 82 16763 134
rect 18950 0 18996 254
rect 19195 82 19201 134
rect 19253 82 19259 134
rect 21446 0 21492 254
rect 21691 82 21697 134
rect 21749 82 21755 134
rect 23942 0 23988 254
rect 24187 82 24193 134
rect 24245 82 24251 134
rect 26438 0 26484 254
rect 26683 82 26689 134
rect 26741 82 26747 134
rect 28934 0 28980 254
rect 29179 82 29185 134
rect 29237 82 29243 134
rect 31430 0 31476 254
rect 31675 82 31681 134
rect 31733 82 31739 134
rect 33926 0 33972 254
rect 34171 82 34177 134
rect 34229 82 34235 134
rect 36422 0 36468 254
rect 36667 82 36673 134
rect 36725 82 36731 134
rect 38918 0 38964 254
rect 39163 82 39169 134
rect 39221 82 39227 134
rect 41414 0 41460 254
rect 41659 82 41665 134
rect 41717 82 41723 134
rect 43910 0 43956 254
rect 44155 82 44161 134
rect 44213 82 44219 134
rect 46406 0 46452 254
rect 46651 82 46657 134
rect 46709 82 46715 134
rect 48902 0 48948 254
rect 49147 82 49153 134
rect 49205 82 49211 134
rect 51398 0 51444 254
rect 51643 82 51649 134
rect 51701 82 51707 134
rect 53894 0 53940 254
rect 54139 82 54145 134
rect 54197 82 54203 134
rect 56390 0 56436 254
rect 56635 82 56641 134
rect 56693 82 56699 134
rect 58886 0 58932 254
rect 59131 82 59137 134
rect 59189 82 59195 134
rect 61382 0 61428 254
rect 61627 82 61633 134
rect 61685 82 61691 134
rect 63878 0 63924 254
rect 64123 82 64129 134
rect 64181 82 64187 134
rect 66374 0 66420 254
rect 66619 82 66625 134
rect 66677 82 66683 134
rect 68870 0 68916 254
rect 69115 82 69121 134
rect 69173 82 69179 134
rect 71366 0 71412 254
rect 71611 82 71617 134
rect 71669 82 71675 134
rect 73862 0 73908 254
rect 74107 82 74113 134
rect 74165 82 74171 134
rect 76358 0 76404 254
rect 76603 82 76609 134
rect 76661 82 76667 134
rect 78854 0 78900 254
rect 79099 82 79105 134
rect 79157 82 79163 134
<< via1 >>
rect 1471 2168 1523 2220
rect 3967 2168 4019 2220
rect 1799 2016 1851 2068
rect 1717 1242 1769 1294
rect 6463 2168 6515 2220
rect 4295 2016 4347 2068
rect 4213 1242 4265 1294
rect 8959 2168 9011 2220
rect 6791 2016 6843 2068
rect 6709 1242 6761 1294
rect 11455 2168 11507 2220
rect 9287 2016 9339 2068
rect 9205 1242 9257 1294
rect 13951 2168 14003 2220
rect 11783 2016 11835 2068
rect 11701 1242 11753 1294
rect 16447 2168 16499 2220
rect 14279 2016 14331 2068
rect 14197 1242 14249 1294
rect 18943 2168 18995 2220
rect 16775 2016 16827 2068
rect 16693 1242 16745 1294
rect 21439 2168 21491 2220
rect 19271 2016 19323 2068
rect 19189 1242 19241 1294
rect 23935 2168 23987 2220
rect 21767 2016 21819 2068
rect 21685 1242 21737 1294
rect 26431 2168 26483 2220
rect 24263 2016 24315 2068
rect 24181 1242 24233 1294
rect 28927 2168 28979 2220
rect 26759 2016 26811 2068
rect 26677 1242 26729 1294
rect 31423 2168 31475 2220
rect 29255 2016 29307 2068
rect 29173 1242 29225 1294
rect 33919 2168 33971 2220
rect 31751 2016 31803 2068
rect 31669 1242 31721 1294
rect 36415 2168 36467 2220
rect 34247 2016 34299 2068
rect 34165 1242 34217 1294
rect 38911 2168 38963 2220
rect 36743 2016 36795 2068
rect 36661 1242 36713 1294
rect 41407 2168 41459 2220
rect 39239 2016 39291 2068
rect 39157 1242 39209 1294
rect 43903 2168 43955 2220
rect 41735 2016 41787 2068
rect 41653 1242 41705 1294
rect 46399 2168 46451 2220
rect 44231 2016 44283 2068
rect 44149 1242 44201 1294
rect 48895 2168 48947 2220
rect 46727 2016 46779 2068
rect 46645 1242 46697 1294
rect 51391 2168 51443 2220
rect 49223 2016 49275 2068
rect 49141 1242 49193 1294
rect 53887 2168 53939 2220
rect 51719 2016 51771 2068
rect 51637 1242 51689 1294
rect 56383 2168 56435 2220
rect 54215 2016 54267 2068
rect 54133 1242 54185 1294
rect 58879 2168 58931 2220
rect 56711 2016 56763 2068
rect 56629 1242 56681 1294
rect 61375 2168 61427 2220
rect 59207 2016 59259 2068
rect 59125 1242 59177 1294
rect 63871 2168 63923 2220
rect 61703 2016 61755 2068
rect 61621 1242 61673 1294
rect 66367 2168 66419 2220
rect 64199 2016 64251 2068
rect 64117 1242 64169 1294
rect 68863 2168 68915 2220
rect 66695 2016 66747 2068
rect 66613 1242 66665 1294
rect 71359 2168 71411 2220
rect 69191 2016 69243 2068
rect 69109 1242 69161 1294
rect 73855 2168 73907 2220
rect 71687 2016 71739 2068
rect 71605 1242 71657 1294
rect 76351 2168 76403 2220
rect 74183 2016 74235 2068
rect 74101 1242 74153 1294
rect 78847 2168 78899 2220
rect 76679 2016 76731 2068
rect 76597 1242 76649 1294
rect 79175 2016 79227 2068
rect 79093 1242 79145 1294
rect 1729 404 1781 456
rect 4225 404 4277 456
rect 6721 404 6773 456
rect 9217 404 9269 456
rect 11713 404 11765 456
rect 14209 404 14261 456
rect 16705 404 16757 456
rect 19201 404 19253 456
rect 21697 404 21749 456
rect 24193 404 24245 456
rect 26689 404 26741 456
rect 29185 404 29237 456
rect 31681 404 31733 456
rect 34177 404 34229 456
rect 36673 404 36725 456
rect 39169 404 39221 456
rect 41665 404 41717 456
rect 44161 404 44213 456
rect 46657 404 46709 456
rect 49153 404 49205 456
rect 51649 404 51701 456
rect 54145 404 54197 456
rect 56641 404 56693 456
rect 59137 404 59189 456
rect 61633 404 61685 456
rect 64129 404 64181 456
rect 66625 404 66677 456
rect 69121 404 69173 456
rect 71617 404 71669 456
rect 74113 404 74165 456
rect 76609 404 76661 456
rect 79105 404 79157 456
rect 1729 82 1781 134
rect 4225 82 4277 134
rect 6721 82 6773 134
rect 9217 82 9269 134
rect 11713 82 11765 134
rect 14209 82 14261 134
rect 16705 82 16757 134
rect 19201 82 19253 134
rect 21697 82 21749 134
rect 24193 82 24245 134
rect 26689 82 26741 134
rect 29185 82 29237 134
rect 31681 82 31733 134
rect 34177 82 34229 134
rect 36673 82 36725 134
rect 39169 82 39221 134
rect 41665 82 41717 134
rect 44161 82 44213 134
rect 46657 82 46709 134
rect 49153 82 49205 134
rect 51649 82 51701 134
rect 54145 82 54197 134
rect 56641 82 56693 134
rect 59137 82 59189 134
rect 61633 82 61685 134
rect 64129 82 64181 134
rect 66625 82 66677 134
rect 69121 82 69173 134
rect 71617 82 71669 134
rect 74113 82 74165 134
rect 76609 82 76661 134
rect 79105 82 79157 134
<< metal2 >>
rect 1469 2222 1525 2231
rect 1469 2157 1525 2166
rect 3965 2222 4021 2231
rect 3965 2157 4021 2166
rect 6461 2222 6517 2231
rect 6461 2157 6517 2166
rect 8957 2222 9013 2231
rect 8957 2157 9013 2166
rect 11453 2222 11509 2231
rect 11453 2157 11509 2166
rect 13949 2222 14005 2231
rect 13949 2157 14005 2166
rect 16445 2222 16501 2231
rect 16445 2157 16501 2166
rect 18941 2222 18997 2231
rect 18941 2157 18997 2166
rect 21437 2222 21493 2231
rect 21437 2157 21493 2166
rect 23933 2222 23989 2231
rect 23933 2157 23989 2166
rect 26429 2222 26485 2231
rect 26429 2157 26485 2166
rect 28925 2222 28981 2231
rect 28925 2157 28981 2166
rect 31421 2222 31477 2231
rect 31421 2157 31477 2166
rect 33917 2222 33973 2231
rect 33917 2157 33973 2166
rect 36413 2222 36469 2231
rect 36413 2157 36469 2166
rect 38909 2222 38965 2231
rect 38909 2157 38965 2166
rect 41405 2222 41461 2231
rect 41405 2157 41461 2166
rect 43901 2222 43957 2231
rect 43901 2157 43957 2166
rect 46397 2222 46453 2231
rect 46397 2157 46453 2166
rect 48893 2222 48949 2231
rect 48893 2157 48949 2166
rect 51389 2222 51445 2231
rect 51389 2157 51445 2166
rect 53885 2222 53941 2231
rect 53885 2157 53941 2166
rect 56381 2222 56437 2231
rect 56381 2157 56437 2166
rect 58877 2222 58933 2231
rect 58877 2157 58933 2166
rect 61373 2222 61429 2231
rect 61373 2157 61429 2166
rect 63869 2222 63925 2231
rect 63869 2157 63925 2166
rect 66365 2222 66421 2231
rect 66365 2157 66421 2166
rect 68861 2222 68917 2231
rect 68861 2157 68917 2166
rect 71357 2222 71413 2231
rect 71357 2157 71413 2166
rect 73853 2222 73909 2231
rect 73853 2157 73909 2166
rect 76349 2222 76405 2231
rect 76349 2157 76405 2166
rect 78845 2222 78901 2231
rect 78845 2157 78901 2166
rect 1797 2070 1853 2079
rect 1797 2005 1853 2014
rect 4293 2070 4349 2079
rect 4293 2005 4349 2014
rect 6789 2070 6845 2079
rect 6789 2005 6845 2014
rect 9285 2070 9341 2079
rect 9285 2005 9341 2014
rect 11781 2070 11837 2079
rect 11781 2005 11837 2014
rect 14277 2070 14333 2079
rect 14277 2005 14333 2014
rect 16773 2070 16829 2079
rect 16773 2005 16829 2014
rect 19269 2070 19325 2079
rect 19269 2005 19325 2014
rect 21765 2070 21821 2079
rect 21765 2005 21821 2014
rect 24261 2070 24317 2079
rect 24261 2005 24317 2014
rect 26757 2070 26813 2079
rect 26757 2005 26813 2014
rect 29253 2070 29309 2079
rect 29253 2005 29309 2014
rect 31749 2070 31805 2079
rect 31749 2005 31805 2014
rect 34245 2070 34301 2079
rect 34245 2005 34301 2014
rect 36741 2070 36797 2079
rect 36741 2005 36797 2014
rect 39237 2070 39293 2079
rect 39237 2005 39293 2014
rect 41733 2070 41789 2079
rect 41733 2005 41789 2014
rect 44229 2070 44285 2079
rect 44229 2005 44285 2014
rect 46725 2070 46781 2079
rect 46725 2005 46781 2014
rect 49221 2070 49277 2079
rect 49221 2005 49277 2014
rect 51717 2070 51773 2079
rect 51717 2005 51773 2014
rect 54213 2070 54269 2079
rect 54213 2005 54269 2014
rect 56709 2070 56765 2079
rect 56709 2005 56765 2014
rect 59205 2070 59261 2079
rect 59205 2005 59261 2014
rect 61701 2070 61757 2079
rect 61701 2005 61757 2014
rect 64197 2070 64253 2079
rect 64197 2005 64253 2014
rect 66693 2070 66749 2079
rect 66693 2005 66749 2014
rect 69189 2070 69245 2079
rect 69189 2005 69245 2014
rect 71685 2070 71741 2079
rect 71685 2005 71741 2014
rect 74181 2070 74237 2079
rect 74181 2005 74237 2014
rect 76677 2070 76733 2079
rect 76677 2005 76733 2014
rect 79173 2070 79229 2079
rect 79173 2005 79229 2014
rect 1715 1296 1771 1305
rect 1715 1231 1771 1240
rect 4211 1296 4267 1305
rect 4211 1231 4267 1240
rect 6707 1296 6763 1305
rect 6707 1231 6763 1240
rect 9203 1296 9259 1305
rect 9203 1231 9259 1240
rect 11699 1296 11755 1305
rect 11699 1231 11755 1240
rect 14195 1296 14251 1305
rect 14195 1231 14251 1240
rect 16691 1296 16747 1305
rect 16691 1231 16747 1240
rect 19187 1296 19243 1305
rect 19187 1231 19243 1240
rect 21683 1296 21739 1305
rect 21683 1231 21739 1240
rect 24179 1296 24235 1305
rect 24179 1231 24235 1240
rect 26675 1296 26731 1305
rect 26675 1231 26731 1240
rect 29171 1296 29227 1305
rect 29171 1231 29227 1240
rect 31667 1296 31723 1305
rect 31667 1231 31723 1240
rect 34163 1296 34219 1305
rect 34163 1231 34219 1240
rect 36659 1296 36715 1305
rect 36659 1231 36715 1240
rect 39155 1296 39211 1305
rect 39155 1231 39211 1240
rect 41651 1296 41707 1305
rect 41651 1231 41707 1240
rect 44147 1296 44203 1305
rect 44147 1231 44203 1240
rect 46643 1296 46699 1305
rect 46643 1231 46699 1240
rect 49139 1296 49195 1305
rect 49139 1231 49195 1240
rect 51635 1296 51691 1305
rect 51635 1231 51691 1240
rect 54131 1296 54187 1305
rect 54131 1231 54187 1240
rect 56627 1296 56683 1305
rect 56627 1231 56683 1240
rect 59123 1296 59179 1305
rect 59123 1231 59179 1240
rect 61619 1296 61675 1305
rect 61619 1231 61675 1240
rect 64115 1296 64171 1305
rect 64115 1231 64171 1240
rect 66611 1296 66667 1305
rect 66611 1231 66667 1240
rect 69107 1296 69163 1305
rect 69107 1231 69163 1240
rect 71603 1296 71659 1305
rect 71603 1231 71659 1240
rect 74099 1296 74155 1305
rect 74099 1231 74155 1240
rect 76595 1296 76651 1305
rect 76595 1231 76651 1240
rect 79091 1296 79147 1305
rect 79091 1231 79147 1240
rect 1727 458 1783 467
rect 1727 393 1783 402
rect 4223 458 4279 467
rect 4223 393 4279 402
rect 6719 458 6775 467
rect 6719 393 6775 402
rect 9215 458 9271 467
rect 9215 393 9271 402
rect 11711 458 11767 467
rect 11711 393 11767 402
rect 14207 458 14263 467
rect 14207 393 14263 402
rect 16703 458 16759 467
rect 16703 393 16759 402
rect 19199 458 19255 467
rect 19199 393 19255 402
rect 21695 458 21751 467
rect 21695 393 21751 402
rect 24191 458 24247 467
rect 24191 393 24247 402
rect 26687 458 26743 467
rect 26687 393 26743 402
rect 29183 458 29239 467
rect 29183 393 29239 402
rect 31679 458 31735 467
rect 31679 393 31735 402
rect 34175 458 34231 467
rect 34175 393 34231 402
rect 36671 458 36727 467
rect 36671 393 36727 402
rect 39167 458 39223 467
rect 39167 393 39223 402
rect 41663 458 41719 467
rect 41663 393 41719 402
rect 44159 458 44215 467
rect 44159 393 44215 402
rect 46655 458 46711 467
rect 46655 393 46711 402
rect 49151 458 49207 467
rect 49151 393 49207 402
rect 51647 458 51703 467
rect 51647 393 51703 402
rect 54143 458 54199 467
rect 54143 393 54199 402
rect 56639 458 56695 467
rect 56639 393 56695 402
rect 59135 458 59191 467
rect 59135 393 59191 402
rect 61631 458 61687 467
rect 61631 393 61687 402
rect 64127 458 64183 467
rect 64127 393 64183 402
rect 66623 458 66679 467
rect 66623 393 66679 402
rect 69119 458 69175 467
rect 69119 393 69175 402
rect 71615 458 71671 467
rect 71615 393 71671 402
rect 74111 458 74167 467
rect 74111 393 74167 402
rect 76607 458 76663 467
rect 76607 393 76663 402
rect 79103 458 79159 467
rect 79103 393 79159 402
rect 1727 136 1783 145
rect 1727 71 1783 80
rect 4223 136 4279 145
rect 4223 71 4279 80
rect 6719 136 6775 145
rect 6719 71 6775 80
rect 9215 136 9271 145
rect 9215 71 9271 80
rect 11711 136 11767 145
rect 11711 71 11767 80
rect 14207 136 14263 145
rect 14207 71 14263 80
rect 16703 136 16759 145
rect 16703 71 16759 80
rect 19199 136 19255 145
rect 19199 71 19255 80
rect 21695 136 21751 145
rect 21695 71 21751 80
rect 24191 136 24247 145
rect 24191 71 24247 80
rect 26687 136 26743 145
rect 26687 71 26743 80
rect 29183 136 29239 145
rect 29183 71 29239 80
rect 31679 136 31735 145
rect 31679 71 31735 80
rect 34175 136 34231 145
rect 34175 71 34231 80
rect 36671 136 36727 145
rect 36671 71 36727 80
rect 39167 136 39223 145
rect 39167 71 39223 80
rect 41663 136 41719 145
rect 41663 71 41719 80
rect 44159 136 44215 145
rect 44159 71 44215 80
rect 46655 136 46711 145
rect 46655 71 46711 80
rect 49151 136 49207 145
rect 49151 71 49207 80
rect 51647 136 51703 145
rect 51647 71 51703 80
rect 54143 136 54199 145
rect 54143 71 54199 80
rect 56639 136 56695 145
rect 56639 71 56695 80
rect 59135 136 59191 145
rect 59135 71 59191 80
rect 61631 136 61687 145
rect 61631 71 61687 80
rect 64127 136 64183 145
rect 64127 71 64183 80
rect 66623 136 66679 145
rect 66623 71 66679 80
rect 69119 136 69175 145
rect 69119 71 69175 80
rect 71615 136 71671 145
rect 71615 71 71671 80
rect 74111 136 74167 145
rect 74111 71 74167 80
rect 76607 136 76663 145
rect 76607 71 76663 80
rect 79103 136 79159 145
rect 79103 71 79159 80
<< via2 >>
rect 1469 2220 1525 2222
rect 1469 2168 1471 2220
rect 1471 2168 1523 2220
rect 1523 2168 1525 2220
rect 1469 2166 1525 2168
rect 3965 2220 4021 2222
rect 3965 2168 3967 2220
rect 3967 2168 4019 2220
rect 4019 2168 4021 2220
rect 3965 2166 4021 2168
rect 6461 2220 6517 2222
rect 6461 2168 6463 2220
rect 6463 2168 6515 2220
rect 6515 2168 6517 2220
rect 6461 2166 6517 2168
rect 8957 2220 9013 2222
rect 8957 2168 8959 2220
rect 8959 2168 9011 2220
rect 9011 2168 9013 2220
rect 8957 2166 9013 2168
rect 11453 2220 11509 2222
rect 11453 2168 11455 2220
rect 11455 2168 11507 2220
rect 11507 2168 11509 2220
rect 11453 2166 11509 2168
rect 13949 2220 14005 2222
rect 13949 2168 13951 2220
rect 13951 2168 14003 2220
rect 14003 2168 14005 2220
rect 13949 2166 14005 2168
rect 16445 2220 16501 2222
rect 16445 2168 16447 2220
rect 16447 2168 16499 2220
rect 16499 2168 16501 2220
rect 16445 2166 16501 2168
rect 18941 2220 18997 2222
rect 18941 2168 18943 2220
rect 18943 2168 18995 2220
rect 18995 2168 18997 2220
rect 18941 2166 18997 2168
rect 21437 2220 21493 2222
rect 21437 2168 21439 2220
rect 21439 2168 21491 2220
rect 21491 2168 21493 2220
rect 21437 2166 21493 2168
rect 23933 2220 23989 2222
rect 23933 2168 23935 2220
rect 23935 2168 23987 2220
rect 23987 2168 23989 2220
rect 23933 2166 23989 2168
rect 26429 2220 26485 2222
rect 26429 2168 26431 2220
rect 26431 2168 26483 2220
rect 26483 2168 26485 2220
rect 26429 2166 26485 2168
rect 28925 2220 28981 2222
rect 28925 2168 28927 2220
rect 28927 2168 28979 2220
rect 28979 2168 28981 2220
rect 28925 2166 28981 2168
rect 31421 2220 31477 2222
rect 31421 2168 31423 2220
rect 31423 2168 31475 2220
rect 31475 2168 31477 2220
rect 31421 2166 31477 2168
rect 33917 2220 33973 2222
rect 33917 2168 33919 2220
rect 33919 2168 33971 2220
rect 33971 2168 33973 2220
rect 33917 2166 33973 2168
rect 36413 2220 36469 2222
rect 36413 2168 36415 2220
rect 36415 2168 36467 2220
rect 36467 2168 36469 2220
rect 36413 2166 36469 2168
rect 38909 2220 38965 2222
rect 38909 2168 38911 2220
rect 38911 2168 38963 2220
rect 38963 2168 38965 2220
rect 38909 2166 38965 2168
rect 41405 2220 41461 2222
rect 41405 2168 41407 2220
rect 41407 2168 41459 2220
rect 41459 2168 41461 2220
rect 41405 2166 41461 2168
rect 43901 2220 43957 2222
rect 43901 2168 43903 2220
rect 43903 2168 43955 2220
rect 43955 2168 43957 2220
rect 43901 2166 43957 2168
rect 46397 2220 46453 2222
rect 46397 2168 46399 2220
rect 46399 2168 46451 2220
rect 46451 2168 46453 2220
rect 46397 2166 46453 2168
rect 48893 2220 48949 2222
rect 48893 2168 48895 2220
rect 48895 2168 48947 2220
rect 48947 2168 48949 2220
rect 48893 2166 48949 2168
rect 51389 2220 51445 2222
rect 51389 2168 51391 2220
rect 51391 2168 51443 2220
rect 51443 2168 51445 2220
rect 51389 2166 51445 2168
rect 53885 2220 53941 2222
rect 53885 2168 53887 2220
rect 53887 2168 53939 2220
rect 53939 2168 53941 2220
rect 53885 2166 53941 2168
rect 56381 2220 56437 2222
rect 56381 2168 56383 2220
rect 56383 2168 56435 2220
rect 56435 2168 56437 2220
rect 56381 2166 56437 2168
rect 58877 2220 58933 2222
rect 58877 2168 58879 2220
rect 58879 2168 58931 2220
rect 58931 2168 58933 2220
rect 58877 2166 58933 2168
rect 61373 2220 61429 2222
rect 61373 2168 61375 2220
rect 61375 2168 61427 2220
rect 61427 2168 61429 2220
rect 61373 2166 61429 2168
rect 63869 2220 63925 2222
rect 63869 2168 63871 2220
rect 63871 2168 63923 2220
rect 63923 2168 63925 2220
rect 63869 2166 63925 2168
rect 66365 2220 66421 2222
rect 66365 2168 66367 2220
rect 66367 2168 66419 2220
rect 66419 2168 66421 2220
rect 66365 2166 66421 2168
rect 68861 2220 68917 2222
rect 68861 2168 68863 2220
rect 68863 2168 68915 2220
rect 68915 2168 68917 2220
rect 68861 2166 68917 2168
rect 71357 2220 71413 2222
rect 71357 2168 71359 2220
rect 71359 2168 71411 2220
rect 71411 2168 71413 2220
rect 71357 2166 71413 2168
rect 73853 2220 73909 2222
rect 73853 2168 73855 2220
rect 73855 2168 73907 2220
rect 73907 2168 73909 2220
rect 73853 2166 73909 2168
rect 76349 2220 76405 2222
rect 76349 2168 76351 2220
rect 76351 2168 76403 2220
rect 76403 2168 76405 2220
rect 76349 2166 76405 2168
rect 78845 2220 78901 2222
rect 78845 2168 78847 2220
rect 78847 2168 78899 2220
rect 78899 2168 78901 2220
rect 78845 2166 78901 2168
rect 1797 2068 1853 2070
rect 1797 2016 1799 2068
rect 1799 2016 1851 2068
rect 1851 2016 1853 2068
rect 1797 2014 1853 2016
rect 4293 2068 4349 2070
rect 4293 2016 4295 2068
rect 4295 2016 4347 2068
rect 4347 2016 4349 2068
rect 4293 2014 4349 2016
rect 6789 2068 6845 2070
rect 6789 2016 6791 2068
rect 6791 2016 6843 2068
rect 6843 2016 6845 2068
rect 6789 2014 6845 2016
rect 9285 2068 9341 2070
rect 9285 2016 9287 2068
rect 9287 2016 9339 2068
rect 9339 2016 9341 2068
rect 9285 2014 9341 2016
rect 11781 2068 11837 2070
rect 11781 2016 11783 2068
rect 11783 2016 11835 2068
rect 11835 2016 11837 2068
rect 11781 2014 11837 2016
rect 14277 2068 14333 2070
rect 14277 2016 14279 2068
rect 14279 2016 14331 2068
rect 14331 2016 14333 2068
rect 14277 2014 14333 2016
rect 16773 2068 16829 2070
rect 16773 2016 16775 2068
rect 16775 2016 16827 2068
rect 16827 2016 16829 2068
rect 16773 2014 16829 2016
rect 19269 2068 19325 2070
rect 19269 2016 19271 2068
rect 19271 2016 19323 2068
rect 19323 2016 19325 2068
rect 19269 2014 19325 2016
rect 21765 2068 21821 2070
rect 21765 2016 21767 2068
rect 21767 2016 21819 2068
rect 21819 2016 21821 2068
rect 21765 2014 21821 2016
rect 24261 2068 24317 2070
rect 24261 2016 24263 2068
rect 24263 2016 24315 2068
rect 24315 2016 24317 2068
rect 24261 2014 24317 2016
rect 26757 2068 26813 2070
rect 26757 2016 26759 2068
rect 26759 2016 26811 2068
rect 26811 2016 26813 2068
rect 26757 2014 26813 2016
rect 29253 2068 29309 2070
rect 29253 2016 29255 2068
rect 29255 2016 29307 2068
rect 29307 2016 29309 2068
rect 29253 2014 29309 2016
rect 31749 2068 31805 2070
rect 31749 2016 31751 2068
rect 31751 2016 31803 2068
rect 31803 2016 31805 2068
rect 31749 2014 31805 2016
rect 34245 2068 34301 2070
rect 34245 2016 34247 2068
rect 34247 2016 34299 2068
rect 34299 2016 34301 2068
rect 34245 2014 34301 2016
rect 36741 2068 36797 2070
rect 36741 2016 36743 2068
rect 36743 2016 36795 2068
rect 36795 2016 36797 2068
rect 36741 2014 36797 2016
rect 39237 2068 39293 2070
rect 39237 2016 39239 2068
rect 39239 2016 39291 2068
rect 39291 2016 39293 2068
rect 39237 2014 39293 2016
rect 41733 2068 41789 2070
rect 41733 2016 41735 2068
rect 41735 2016 41787 2068
rect 41787 2016 41789 2068
rect 41733 2014 41789 2016
rect 44229 2068 44285 2070
rect 44229 2016 44231 2068
rect 44231 2016 44283 2068
rect 44283 2016 44285 2068
rect 44229 2014 44285 2016
rect 46725 2068 46781 2070
rect 46725 2016 46727 2068
rect 46727 2016 46779 2068
rect 46779 2016 46781 2068
rect 46725 2014 46781 2016
rect 49221 2068 49277 2070
rect 49221 2016 49223 2068
rect 49223 2016 49275 2068
rect 49275 2016 49277 2068
rect 49221 2014 49277 2016
rect 51717 2068 51773 2070
rect 51717 2016 51719 2068
rect 51719 2016 51771 2068
rect 51771 2016 51773 2068
rect 51717 2014 51773 2016
rect 54213 2068 54269 2070
rect 54213 2016 54215 2068
rect 54215 2016 54267 2068
rect 54267 2016 54269 2068
rect 54213 2014 54269 2016
rect 56709 2068 56765 2070
rect 56709 2016 56711 2068
rect 56711 2016 56763 2068
rect 56763 2016 56765 2068
rect 56709 2014 56765 2016
rect 59205 2068 59261 2070
rect 59205 2016 59207 2068
rect 59207 2016 59259 2068
rect 59259 2016 59261 2068
rect 59205 2014 59261 2016
rect 61701 2068 61757 2070
rect 61701 2016 61703 2068
rect 61703 2016 61755 2068
rect 61755 2016 61757 2068
rect 61701 2014 61757 2016
rect 64197 2068 64253 2070
rect 64197 2016 64199 2068
rect 64199 2016 64251 2068
rect 64251 2016 64253 2068
rect 64197 2014 64253 2016
rect 66693 2068 66749 2070
rect 66693 2016 66695 2068
rect 66695 2016 66747 2068
rect 66747 2016 66749 2068
rect 66693 2014 66749 2016
rect 69189 2068 69245 2070
rect 69189 2016 69191 2068
rect 69191 2016 69243 2068
rect 69243 2016 69245 2068
rect 69189 2014 69245 2016
rect 71685 2068 71741 2070
rect 71685 2016 71687 2068
rect 71687 2016 71739 2068
rect 71739 2016 71741 2068
rect 71685 2014 71741 2016
rect 74181 2068 74237 2070
rect 74181 2016 74183 2068
rect 74183 2016 74235 2068
rect 74235 2016 74237 2068
rect 74181 2014 74237 2016
rect 76677 2068 76733 2070
rect 76677 2016 76679 2068
rect 76679 2016 76731 2068
rect 76731 2016 76733 2068
rect 76677 2014 76733 2016
rect 79173 2068 79229 2070
rect 79173 2016 79175 2068
rect 79175 2016 79227 2068
rect 79227 2016 79229 2068
rect 79173 2014 79229 2016
rect 1715 1294 1771 1296
rect 1715 1242 1717 1294
rect 1717 1242 1769 1294
rect 1769 1242 1771 1294
rect 1715 1240 1771 1242
rect 4211 1294 4267 1296
rect 4211 1242 4213 1294
rect 4213 1242 4265 1294
rect 4265 1242 4267 1294
rect 4211 1240 4267 1242
rect 6707 1294 6763 1296
rect 6707 1242 6709 1294
rect 6709 1242 6761 1294
rect 6761 1242 6763 1294
rect 6707 1240 6763 1242
rect 9203 1294 9259 1296
rect 9203 1242 9205 1294
rect 9205 1242 9257 1294
rect 9257 1242 9259 1294
rect 9203 1240 9259 1242
rect 11699 1294 11755 1296
rect 11699 1242 11701 1294
rect 11701 1242 11753 1294
rect 11753 1242 11755 1294
rect 11699 1240 11755 1242
rect 14195 1294 14251 1296
rect 14195 1242 14197 1294
rect 14197 1242 14249 1294
rect 14249 1242 14251 1294
rect 14195 1240 14251 1242
rect 16691 1294 16747 1296
rect 16691 1242 16693 1294
rect 16693 1242 16745 1294
rect 16745 1242 16747 1294
rect 16691 1240 16747 1242
rect 19187 1294 19243 1296
rect 19187 1242 19189 1294
rect 19189 1242 19241 1294
rect 19241 1242 19243 1294
rect 19187 1240 19243 1242
rect 21683 1294 21739 1296
rect 21683 1242 21685 1294
rect 21685 1242 21737 1294
rect 21737 1242 21739 1294
rect 21683 1240 21739 1242
rect 24179 1294 24235 1296
rect 24179 1242 24181 1294
rect 24181 1242 24233 1294
rect 24233 1242 24235 1294
rect 24179 1240 24235 1242
rect 26675 1294 26731 1296
rect 26675 1242 26677 1294
rect 26677 1242 26729 1294
rect 26729 1242 26731 1294
rect 26675 1240 26731 1242
rect 29171 1294 29227 1296
rect 29171 1242 29173 1294
rect 29173 1242 29225 1294
rect 29225 1242 29227 1294
rect 29171 1240 29227 1242
rect 31667 1294 31723 1296
rect 31667 1242 31669 1294
rect 31669 1242 31721 1294
rect 31721 1242 31723 1294
rect 31667 1240 31723 1242
rect 34163 1294 34219 1296
rect 34163 1242 34165 1294
rect 34165 1242 34217 1294
rect 34217 1242 34219 1294
rect 34163 1240 34219 1242
rect 36659 1294 36715 1296
rect 36659 1242 36661 1294
rect 36661 1242 36713 1294
rect 36713 1242 36715 1294
rect 36659 1240 36715 1242
rect 39155 1294 39211 1296
rect 39155 1242 39157 1294
rect 39157 1242 39209 1294
rect 39209 1242 39211 1294
rect 39155 1240 39211 1242
rect 41651 1294 41707 1296
rect 41651 1242 41653 1294
rect 41653 1242 41705 1294
rect 41705 1242 41707 1294
rect 41651 1240 41707 1242
rect 44147 1294 44203 1296
rect 44147 1242 44149 1294
rect 44149 1242 44201 1294
rect 44201 1242 44203 1294
rect 44147 1240 44203 1242
rect 46643 1294 46699 1296
rect 46643 1242 46645 1294
rect 46645 1242 46697 1294
rect 46697 1242 46699 1294
rect 46643 1240 46699 1242
rect 49139 1294 49195 1296
rect 49139 1242 49141 1294
rect 49141 1242 49193 1294
rect 49193 1242 49195 1294
rect 49139 1240 49195 1242
rect 51635 1294 51691 1296
rect 51635 1242 51637 1294
rect 51637 1242 51689 1294
rect 51689 1242 51691 1294
rect 51635 1240 51691 1242
rect 54131 1294 54187 1296
rect 54131 1242 54133 1294
rect 54133 1242 54185 1294
rect 54185 1242 54187 1294
rect 54131 1240 54187 1242
rect 56627 1294 56683 1296
rect 56627 1242 56629 1294
rect 56629 1242 56681 1294
rect 56681 1242 56683 1294
rect 56627 1240 56683 1242
rect 59123 1294 59179 1296
rect 59123 1242 59125 1294
rect 59125 1242 59177 1294
rect 59177 1242 59179 1294
rect 59123 1240 59179 1242
rect 61619 1294 61675 1296
rect 61619 1242 61621 1294
rect 61621 1242 61673 1294
rect 61673 1242 61675 1294
rect 61619 1240 61675 1242
rect 64115 1294 64171 1296
rect 64115 1242 64117 1294
rect 64117 1242 64169 1294
rect 64169 1242 64171 1294
rect 64115 1240 64171 1242
rect 66611 1294 66667 1296
rect 66611 1242 66613 1294
rect 66613 1242 66665 1294
rect 66665 1242 66667 1294
rect 66611 1240 66667 1242
rect 69107 1294 69163 1296
rect 69107 1242 69109 1294
rect 69109 1242 69161 1294
rect 69161 1242 69163 1294
rect 69107 1240 69163 1242
rect 71603 1294 71659 1296
rect 71603 1242 71605 1294
rect 71605 1242 71657 1294
rect 71657 1242 71659 1294
rect 71603 1240 71659 1242
rect 74099 1294 74155 1296
rect 74099 1242 74101 1294
rect 74101 1242 74153 1294
rect 74153 1242 74155 1294
rect 74099 1240 74155 1242
rect 76595 1294 76651 1296
rect 76595 1242 76597 1294
rect 76597 1242 76649 1294
rect 76649 1242 76651 1294
rect 76595 1240 76651 1242
rect 79091 1294 79147 1296
rect 79091 1242 79093 1294
rect 79093 1242 79145 1294
rect 79145 1242 79147 1294
rect 79091 1240 79147 1242
rect 1727 456 1783 458
rect 1727 404 1729 456
rect 1729 404 1781 456
rect 1781 404 1783 456
rect 1727 402 1783 404
rect 4223 456 4279 458
rect 4223 404 4225 456
rect 4225 404 4277 456
rect 4277 404 4279 456
rect 4223 402 4279 404
rect 6719 456 6775 458
rect 6719 404 6721 456
rect 6721 404 6773 456
rect 6773 404 6775 456
rect 6719 402 6775 404
rect 9215 456 9271 458
rect 9215 404 9217 456
rect 9217 404 9269 456
rect 9269 404 9271 456
rect 9215 402 9271 404
rect 11711 456 11767 458
rect 11711 404 11713 456
rect 11713 404 11765 456
rect 11765 404 11767 456
rect 11711 402 11767 404
rect 14207 456 14263 458
rect 14207 404 14209 456
rect 14209 404 14261 456
rect 14261 404 14263 456
rect 14207 402 14263 404
rect 16703 456 16759 458
rect 16703 404 16705 456
rect 16705 404 16757 456
rect 16757 404 16759 456
rect 16703 402 16759 404
rect 19199 456 19255 458
rect 19199 404 19201 456
rect 19201 404 19253 456
rect 19253 404 19255 456
rect 19199 402 19255 404
rect 21695 456 21751 458
rect 21695 404 21697 456
rect 21697 404 21749 456
rect 21749 404 21751 456
rect 21695 402 21751 404
rect 24191 456 24247 458
rect 24191 404 24193 456
rect 24193 404 24245 456
rect 24245 404 24247 456
rect 24191 402 24247 404
rect 26687 456 26743 458
rect 26687 404 26689 456
rect 26689 404 26741 456
rect 26741 404 26743 456
rect 26687 402 26743 404
rect 29183 456 29239 458
rect 29183 404 29185 456
rect 29185 404 29237 456
rect 29237 404 29239 456
rect 29183 402 29239 404
rect 31679 456 31735 458
rect 31679 404 31681 456
rect 31681 404 31733 456
rect 31733 404 31735 456
rect 31679 402 31735 404
rect 34175 456 34231 458
rect 34175 404 34177 456
rect 34177 404 34229 456
rect 34229 404 34231 456
rect 34175 402 34231 404
rect 36671 456 36727 458
rect 36671 404 36673 456
rect 36673 404 36725 456
rect 36725 404 36727 456
rect 36671 402 36727 404
rect 39167 456 39223 458
rect 39167 404 39169 456
rect 39169 404 39221 456
rect 39221 404 39223 456
rect 39167 402 39223 404
rect 41663 456 41719 458
rect 41663 404 41665 456
rect 41665 404 41717 456
rect 41717 404 41719 456
rect 41663 402 41719 404
rect 44159 456 44215 458
rect 44159 404 44161 456
rect 44161 404 44213 456
rect 44213 404 44215 456
rect 44159 402 44215 404
rect 46655 456 46711 458
rect 46655 404 46657 456
rect 46657 404 46709 456
rect 46709 404 46711 456
rect 46655 402 46711 404
rect 49151 456 49207 458
rect 49151 404 49153 456
rect 49153 404 49205 456
rect 49205 404 49207 456
rect 49151 402 49207 404
rect 51647 456 51703 458
rect 51647 404 51649 456
rect 51649 404 51701 456
rect 51701 404 51703 456
rect 51647 402 51703 404
rect 54143 456 54199 458
rect 54143 404 54145 456
rect 54145 404 54197 456
rect 54197 404 54199 456
rect 54143 402 54199 404
rect 56639 456 56695 458
rect 56639 404 56641 456
rect 56641 404 56693 456
rect 56693 404 56695 456
rect 56639 402 56695 404
rect 59135 456 59191 458
rect 59135 404 59137 456
rect 59137 404 59189 456
rect 59189 404 59191 456
rect 59135 402 59191 404
rect 61631 456 61687 458
rect 61631 404 61633 456
rect 61633 404 61685 456
rect 61685 404 61687 456
rect 61631 402 61687 404
rect 64127 456 64183 458
rect 64127 404 64129 456
rect 64129 404 64181 456
rect 64181 404 64183 456
rect 64127 402 64183 404
rect 66623 456 66679 458
rect 66623 404 66625 456
rect 66625 404 66677 456
rect 66677 404 66679 456
rect 66623 402 66679 404
rect 69119 456 69175 458
rect 69119 404 69121 456
rect 69121 404 69173 456
rect 69173 404 69175 456
rect 69119 402 69175 404
rect 71615 456 71671 458
rect 71615 404 71617 456
rect 71617 404 71669 456
rect 71669 404 71671 456
rect 71615 402 71671 404
rect 74111 456 74167 458
rect 74111 404 74113 456
rect 74113 404 74165 456
rect 74165 404 74167 456
rect 74111 402 74167 404
rect 76607 456 76663 458
rect 76607 404 76609 456
rect 76609 404 76661 456
rect 76661 404 76663 456
rect 76607 402 76663 404
rect 79103 456 79159 458
rect 79103 404 79105 456
rect 79105 404 79157 456
rect 79157 404 79159 456
rect 79103 402 79159 404
rect 1727 134 1783 136
rect 1727 82 1729 134
rect 1729 82 1781 134
rect 1781 82 1783 134
rect 1727 80 1783 82
rect 4223 134 4279 136
rect 4223 82 4225 134
rect 4225 82 4277 134
rect 4277 82 4279 134
rect 4223 80 4279 82
rect 6719 134 6775 136
rect 6719 82 6721 134
rect 6721 82 6773 134
rect 6773 82 6775 134
rect 6719 80 6775 82
rect 9215 134 9271 136
rect 9215 82 9217 134
rect 9217 82 9269 134
rect 9269 82 9271 134
rect 9215 80 9271 82
rect 11711 134 11767 136
rect 11711 82 11713 134
rect 11713 82 11765 134
rect 11765 82 11767 134
rect 11711 80 11767 82
rect 14207 134 14263 136
rect 14207 82 14209 134
rect 14209 82 14261 134
rect 14261 82 14263 134
rect 14207 80 14263 82
rect 16703 134 16759 136
rect 16703 82 16705 134
rect 16705 82 16757 134
rect 16757 82 16759 134
rect 16703 80 16759 82
rect 19199 134 19255 136
rect 19199 82 19201 134
rect 19201 82 19253 134
rect 19253 82 19255 134
rect 19199 80 19255 82
rect 21695 134 21751 136
rect 21695 82 21697 134
rect 21697 82 21749 134
rect 21749 82 21751 134
rect 21695 80 21751 82
rect 24191 134 24247 136
rect 24191 82 24193 134
rect 24193 82 24245 134
rect 24245 82 24247 134
rect 24191 80 24247 82
rect 26687 134 26743 136
rect 26687 82 26689 134
rect 26689 82 26741 134
rect 26741 82 26743 134
rect 26687 80 26743 82
rect 29183 134 29239 136
rect 29183 82 29185 134
rect 29185 82 29237 134
rect 29237 82 29239 134
rect 29183 80 29239 82
rect 31679 134 31735 136
rect 31679 82 31681 134
rect 31681 82 31733 134
rect 31733 82 31735 134
rect 31679 80 31735 82
rect 34175 134 34231 136
rect 34175 82 34177 134
rect 34177 82 34229 134
rect 34229 82 34231 134
rect 34175 80 34231 82
rect 36671 134 36727 136
rect 36671 82 36673 134
rect 36673 82 36725 134
rect 36725 82 36727 134
rect 36671 80 36727 82
rect 39167 134 39223 136
rect 39167 82 39169 134
rect 39169 82 39221 134
rect 39221 82 39223 134
rect 39167 80 39223 82
rect 41663 134 41719 136
rect 41663 82 41665 134
rect 41665 82 41717 134
rect 41717 82 41719 134
rect 41663 80 41719 82
rect 44159 134 44215 136
rect 44159 82 44161 134
rect 44161 82 44213 134
rect 44213 82 44215 134
rect 44159 80 44215 82
rect 46655 134 46711 136
rect 46655 82 46657 134
rect 46657 82 46709 134
rect 46709 82 46711 134
rect 46655 80 46711 82
rect 49151 134 49207 136
rect 49151 82 49153 134
rect 49153 82 49205 134
rect 49205 82 49207 134
rect 49151 80 49207 82
rect 51647 134 51703 136
rect 51647 82 51649 134
rect 51649 82 51701 134
rect 51701 82 51703 134
rect 51647 80 51703 82
rect 54143 134 54199 136
rect 54143 82 54145 134
rect 54145 82 54197 134
rect 54197 82 54199 134
rect 54143 80 54199 82
rect 56639 134 56695 136
rect 56639 82 56641 134
rect 56641 82 56693 134
rect 56693 82 56695 134
rect 56639 80 56695 82
rect 59135 134 59191 136
rect 59135 82 59137 134
rect 59137 82 59189 134
rect 59189 82 59191 134
rect 59135 80 59191 82
rect 61631 134 61687 136
rect 61631 82 61633 134
rect 61633 82 61685 134
rect 61685 82 61687 134
rect 61631 80 61687 82
rect 64127 134 64183 136
rect 64127 82 64129 134
rect 64129 82 64181 134
rect 64181 82 64183 134
rect 64127 80 64183 82
rect 66623 134 66679 136
rect 66623 82 66625 134
rect 66625 82 66677 134
rect 66677 82 66679 134
rect 66623 80 66679 82
rect 69119 134 69175 136
rect 69119 82 69121 134
rect 69121 82 69173 134
rect 69173 82 69175 134
rect 69119 80 69175 82
rect 71615 134 71671 136
rect 71615 82 71617 134
rect 71617 82 71669 134
rect 71669 82 71671 134
rect 71615 80 71671 82
rect 74111 134 74167 136
rect 74111 82 74113 134
rect 74113 82 74165 134
rect 74165 82 74167 134
rect 74111 80 74167 82
rect 76607 134 76663 136
rect 76607 82 76609 134
rect 76609 82 76661 134
rect 76661 82 76663 134
rect 76607 80 76663 82
rect 79103 134 79159 136
rect 79103 82 79105 134
rect 79105 82 79157 134
rect 79157 82 79159 134
rect 79103 80 79159 82
<< metal3 >>
rect 1464 2224 1530 2227
rect 3960 2224 4026 2227
rect 6456 2224 6522 2227
rect 8952 2224 9018 2227
rect 11448 2224 11514 2227
rect 13944 2224 14010 2227
rect 16440 2224 16506 2227
rect 18936 2224 19002 2227
rect 21432 2224 21498 2227
rect 23928 2224 23994 2227
rect 26424 2224 26490 2227
rect 28920 2224 28986 2227
rect 31416 2224 31482 2227
rect 33912 2224 33978 2227
rect 36408 2224 36474 2227
rect 38904 2224 38970 2227
rect 41400 2224 41466 2227
rect 43896 2224 43962 2227
rect 46392 2224 46458 2227
rect 48888 2224 48954 2227
rect 51384 2224 51450 2227
rect 53880 2224 53946 2227
rect 56376 2224 56442 2227
rect 58872 2224 58938 2227
rect 61368 2224 61434 2227
rect 63864 2224 63930 2227
rect 66360 2224 66426 2227
rect 68856 2224 68922 2227
rect 71352 2224 71418 2227
rect 73848 2224 73914 2227
rect 76344 2224 76410 2227
rect 78840 2224 78906 2227
rect 0 2222 79250 2224
rect 0 2166 1469 2222
rect 1525 2166 3965 2222
rect 4021 2166 6461 2222
rect 6517 2166 8957 2222
rect 9013 2166 11453 2222
rect 11509 2166 13949 2222
rect 14005 2166 16445 2222
rect 16501 2166 18941 2222
rect 18997 2166 21437 2222
rect 21493 2166 23933 2222
rect 23989 2166 26429 2222
rect 26485 2166 28925 2222
rect 28981 2166 31421 2222
rect 31477 2166 33917 2222
rect 33973 2166 36413 2222
rect 36469 2166 38909 2222
rect 38965 2166 41405 2222
rect 41461 2166 43901 2222
rect 43957 2166 46397 2222
rect 46453 2166 48893 2222
rect 48949 2166 51389 2222
rect 51445 2166 53885 2222
rect 53941 2166 56381 2222
rect 56437 2166 58877 2222
rect 58933 2166 61373 2222
rect 61429 2166 63869 2222
rect 63925 2166 66365 2222
rect 66421 2166 68861 2222
rect 68917 2166 71357 2222
rect 71413 2166 73853 2222
rect 73909 2166 76349 2222
rect 76405 2166 78845 2222
rect 78901 2166 79250 2222
rect 0 2164 79250 2166
rect 1464 2161 1530 2164
rect 3960 2161 4026 2164
rect 6456 2161 6522 2164
rect 8952 2161 9018 2164
rect 11448 2161 11514 2164
rect 13944 2161 14010 2164
rect 16440 2161 16506 2164
rect 18936 2161 19002 2164
rect 21432 2161 21498 2164
rect 23928 2161 23994 2164
rect 26424 2161 26490 2164
rect 28920 2161 28986 2164
rect 31416 2161 31482 2164
rect 33912 2161 33978 2164
rect 36408 2161 36474 2164
rect 38904 2161 38970 2164
rect 41400 2161 41466 2164
rect 43896 2161 43962 2164
rect 46392 2161 46458 2164
rect 48888 2161 48954 2164
rect 51384 2161 51450 2164
rect 53880 2161 53946 2164
rect 56376 2161 56442 2164
rect 58872 2161 58938 2164
rect 61368 2161 61434 2164
rect 63864 2161 63930 2164
rect 66360 2161 66426 2164
rect 68856 2161 68922 2164
rect 71352 2161 71418 2164
rect 73848 2161 73914 2164
rect 76344 2161 76410 2164
rect 78840 2161 78906 2164
rect 1776 2070 1874 2091
rect 1776 2014 1797 2070
rect 1853 2014 1874 2070
rect 1776 1993 1874 2014
rect 4272 2070 4370 2091
rect 4272 2014 4293 2070
rect 4349 2014 4370 2070
rect 4272 1993 4370 2014
rect 6768 2070 6866 2091
rect 6768 2014 6789 2070
rect 6845 2014 6866 2070
rect 6768 1993 6866 2014
rect 9264 2070 9362 2091
rect 9264 2014 9285 2070
rect 9341 2014 9362 2070
rect 9264 1993 9362 2014
rect 11760 2070 11858 2091
rect 11760 2014 11781 2070
rect 11837 2014 11858 2070
rect 11760 1993 11858 2014
rect 14256 2070 14354 2091
rect 14256 2014 14277 2070
rect 14333 2014 14354 2070
rect 14256 1993 14354 2014
rect 16752 2070 16850 2091
rect 16752 2014 16773 2070
rect 16829 2014 16850 2070
rect 16752 1993 16850 2014
rect 19248 2070 19346 2091
rect 19248 2014 19269 2070
rect 19325 2014 19346 2070
rect 19248 1993 19346 2014
rect 21744 2070 21842 2091
rect 21744 2014 21765 2070
rect 21821 2014 21842 2070
rect 21744 1993 21842 2014
rect 24240 2070 24338 2091
rect 24240 2014 24261 2070
rect 24317 2014 24338 2070
rect 24240 1993 24338 2014
rect 26736 2070 26834 2091
rect 26736 2014 26757 2070
rect 26813 2014 26834 2070
rect 26736 1993 26834 2014
rect 29232 2070 29330 2091
rect 29232 2014 29253 2070
rect 29309 2014 29330 2070
rect 29232 1993 29330 2014
rect 31728 2070 31826 2091
rect 31728 2014 31749 2070
rect 31805 2014 31826 2070
rect 31728 1993 31826 2014
rect 34224 2070 34322 2091
rect 34224 2014 34245 2070
rect 34301 2014 34322 2070
rect 34224 1993 34322 2014
rect 36720 2070 36818 2091
rect 36720 2014 36741 2070
rect 36797 2014 36818 2070
rect 36720 1993 36818 2014
rect 39216 2070 39314 2091
rect 39216 2014 39237 2070
rect 39293 2014 39314 2070
rect 39216 1993 39314 2014
rect 41712 2070 41810 2091
rect 41712 2014 41733 2070
rect 41789 2014 41810 2070
rect 41712 1993 41810 2014
rect 44208 2070 44306 2091
rect 44208 2014 44229 2070
rect 44285 2014 44306 2070
rect 44208 1993 44306 2014
rect 46704 2070 46802 2091
rect 46704 2014 46725 2070
rect 46781 2014 46802 2070
rect 46704 1993 46802 2014
rect 49200 2070 49298 2091
rect 49200 2014 49221 2070
rect 49277 2014 49298 2070
rect 49200 1993 49298 2014
rect 51696 2070 51794 2091
rect 51696 2014 51717 2070
rect 51773 2014 51794 2070
rect 51696 1993 51794 2014
rect 54192 2070 54290 2091
rect 54192 2014 54213 2070
rect 54269 2014 54290 2070
rect 54192 1993 54290 2014
rect 56688 2070 56786 2091
rect 56688 2014 56709 2070
rect 56765 2014 56786 2070
rect 56688 1993 56786 2014
rect 59184 2070 59282 2091
rect 59184 2014 59205 2070
rect 59261 2014 59282 2070
rect 59184 1993 59282 2014
rect 61680 2070 61778 2091
rect 61680 2014 61701 2070
rect 61757 2014 61778 2070
rect 61680 1993 61778 2014
rect 64176 2070 64274 2091
rect 64176 2014 64197 2070
rect 64253 2014 64274 2070
rect 64176 1993 64274 2014
rect 66672 2070 66770 2091
rect 66672 2014 66693 2070
rect 66749 2014 66770 2070
rect 66672 1993 66770 2014
rect 69168 2070 69266 2091
rect 69168 2014 69189 2070
rect 69245 2014 69266 2070
rect 69168 1993 69266 2014
rect 71664 2070 71762 2091
rect 71664 2014 71685 2070
rect 71741 2014 71762 2070
rect 71664 1993 71762 2014
rect 74160 2070 74258 2091
rect 74160 2014 74181 2070
rect 74237 2014 74258 2070
rect 74160 1993 74258 2014
rect 76656 2070 76754 2091
rect 76656 2014 76677 2070
rect 76733 2014 76754 2070
rect 76656 1993 76754 2014
rect 79152 2070 79250 2091
rect 79152 2014 79173 2070
rect 79229 2014 79250 2070
rect 79152 1993 79250 2014
rect 1694 1296 1792 1317
rect 1694 1240 1715 1296
rect 1771 1240 1792 1296
rect 1694 1219 1792 1240
rect 4190 1296 4288 1317
rect 4190 1240 4211 1296
rect 4267 1240 4288 1296
rect 4190 1219 4288 1240
rect 6686 1296 6784 1317
rect 6686 1240 6707 1296
rect 6763 1240 6784 1296
rect 6686 1219 6784 1240
rect 9182 1296 9280 1317
rect 9182 1240 9203 1296
rect 9259 1240 9280 1296
rect 9182 1219 9280 1240
rect 11678 1296 11776 1317
rect 11678 1240 11699 1296
rect 11755 1240 11776 1296
rect 11678 1219 11776 1240
rect 14174 1296 14272 1317
rect 14174 1240 14195 1296
rect 14251 1240 14272 1296
rect 14174 1219 14272 1240
rect 16670 1296 16768 1317
rect 16670 1240 16691 1296
rect 16747 1240 16768 1296
rect 16670 1219 16768 1240
rect 19166 1296 19264 1317
rect 19166 1240 19187 1296
rect 19243 1240 19264 1296
rect 19166 1219 19264 1240
rect 21662 1296 21760 1317
rect 21662 1240 21683 1296
rect 21739 1240 21760 1296
rect 21662 1219 21760 1240
rect 24158 1296 24256 1317
rect 24158 1240 24179 1296
rect 24235 1240 24256 1296
rect 24158 1219 24256 1240
rect 26654 1296 26752 1317
rect 26654 1240 26675 1296
rect 26731 1240 26752 1296
rect 26654 1219 26752 1240
rect 29150 1296 29248 1317
rect 29150 1240 29171 1296
rect 29227 1240 29248 1296
rect 29150 1219 29248 1240
rect 31646 1296 31744 1317
rect 31646 1240 31667 1296
rect 31723 1240 31744 1296
rect 31646 1219 31744 1240
rect 34142 1296 34240 1317
rect 34142 1240 34163 1296
rect 34219 1240 34240 1296
rect 34142 1219 34240 1240
rect 36638 1296 36736 1317
rect 36638 1240 36659 1296
rect 36715 1240 36736 1296
rect 36638 1219 36736 1240
rect 39134 1296 39232 1317
rect 39134 1240 39155 1296
rect 39211 1240 39232 1296
rect 39134 1219 39232 1240
rect 41630 1296 41728 1317
rect 41630 1240 41651 1296
rect 41707 1240 41728 1296
rect 41630 1219 41728 1240
rect 44126 1296 44224 1317
rect 44126 1240 44147 1296
rect 44203 1240 44224 1296
rect 44126 1219 44224 1240
rect 46622 1296 46720 1317
rect 46622 1240 46643 1296
rect 46699 1240 46720 1296
rect 46622 1219 46720 1240
rect 49118 1296 49216 1317
rect 49118 1240 49139 1296
rect 49195 1240 49216 1296
rect 49118 1219 49216 1240
rect 51614 1296 51712 1317
rect 51614 1240 51635 1296
rect 51691 1240 51712 1296
rect 51614 1219 51712 1240
rect 54110 1296 54208 1317
rect 54110 1240 54131 1296
rect 54187 1240 54208 1296
rect 54110 1219 54208 1240
rect 56606 1296 56704 1317
rect 56606 1240 56627 1296
rect 56683 1240 56704 1296
rect 56606 1219 56704 1240
rect 59102 1296 59200 1317
rect 59102 1240 59123 1296
rect 59179 1240 59200 1296
rect 59102 1219 59200 1240
rect 61598 1296 61696 1317
rect 61598 1240 61619 1296
rect 61675 1240 61696 1296
rect 61598 1219 61696 1240
rect 64094 1296 64192 1317
rect 64094 1240 64115 1296
rect 64171 1240 64192 1296
rect 64094 1219 64192 1240
rect 66590 1296 66688 1317
rect 66590 1240 66611 1296
rect 66667 1240 66688 1296
rect 66590 1219 66688 1240
rect 69086 1296 69184 1317
rect 69086 1240 69107 1296
rect 69163 1240 69184 1296
rect 69086 1219 69184 1240
rect 71582 1296 71680 1317
rect 71582 1240 71603 1296
rect 71659 1240 71680 1296
rect 71582 1219 71680 1240
rect 74078 1296 74176 1317
rect 74078 1240 74099 1296
rect 74155 1240 74176 1296
rect 74078 1219 74176 1240
rect 76574 1296 76672 1317
rect 76574 1240 76595 1296
rect 76651 1240 76672 1296
rect 76574 1219 76672 1240
rect 79070 1296 79168 1317
rect 79070 1240 79091 1296
rect 79147 1240 79168 1296
rect 79070 1219 79168 1240
rect 1706 458 1804 479
rect 1706 402 1727 458
rect 1783 402 1804 458
rect 1706 381 1804 402
rect 4202 458 4300 479
rect 4202 402 4223 458
rect 4279 402 4300 458
rect 4202 381 4300 402
rect 6698 458 6796 479
rect 6698 402 6719 458
rect 6775 402 6796 458
rect 6698 381 6796 402
rect 9194 458 9292 479
rect 9194 402 9215 458
rect 9271 402 9292 458
rect 9194 381 9292 402
rect 11690 458 11788 479
rect 11690 402 11711 458
rect 11767 402 11788 458
rect 11690 381 11788 402
rect 14186 458 14284 479
rect 14186 402 14207 458
rect 14263 402 14284 458
rect 14186 381 14284 402
rect 16682 458 16780 479
rect 16682 402 16703 458
rect 16759 402 16780 458
rect 16682 381 16780 402
rect 19178 458 19276 479
rect 19178 402 19199 458
rect 19255 402 19276 458
rect 19178 381 19276 402
rect 21674 458 21772 479
rect 21674 402 21695 458
rect 21751 402 21772 458
rect 21674 381 21772 402
rect 24170 458 24268 479
rect 24170 402 24191 458
rect 24247 402 24268 458
rect 24170 381 24268 402
rect 26666 458 26764 479
rect 26666 402 26687 458
rect 26743 402 26764 458
rect 26666 381 26764 402
rect 29162 458 29260 479
rect 29162 402 29183 458
rect 29239 402 29260 458
rect 29162 381 29260 402
rect 31658 458 31756 479
rect 31658 402 31679 458
rect 31735 402 31756 458
rect 31658 381 31756 402
rect 34154 458 34252 479
rect 34154 402 34175 458
rect 34231 402 34252 458
rect 34154 381 34252 402
rect 36650 458 36748 479
rect 36650 402 36671 458
rect 36727 402 36748 458
rect 36650 381 36748 402
rect 39146 458 39244 479
rect 39146 402 39167 458
rect 39223 402 39244 458
rect 39146 381 39244 402
rect 41642 458 41740 479
rect 41642 402 41663 458
rect 41719 402 41740 458
rect 41642 381 41740 402
rect 44138 458 44236 479
rect 44138 402 44159 458
rect 44215 402 44236 458
rect 44138 381 44236 402
rect 46634 458 46732 479
rect 46634 402 46655 458
rect 46711 402 46732 458
rect 46634 381 46732 402
rect 49130 458 49228 479
rect 49130 402 49151 458
rect 49207 402 49228 458
rect 49130 381 49228 402
rect 51626 458 51724 479
rect 51626 402 51647 458
rect 51703 402 51724 458
rect 51626 381 51724 402
rect 54122 458 54220 479
rect 54122 402 54143 458
rect 54199 402 54220 458
rect 54122 381 54220 402
rect 56618 458 56716 479
rect 56618 402 56639 458
rect 56695 402 56716 458
rect 56618 381 56716 402
rect 59114 458 59212 479
rect 59114 402 59135 458
rect 59191 402 59212 458
rect 59114 381 59212 402
rect 61610 458 61708 479
rect 61610 402 61631 458
rect 61687 402 61708 458
rect 61610 381 61708 402
rect 64106 458 64204 479
rect 64106 402 64127 458
rect 64183 402 64204 458
rect 64106 381 64204 402
rect 66602 458 66700 479
rect 66602 402 66623 458
rect 66679 402 66700 458
rect 66602 381 66700 402
rect 69098 458 69196 479
rect 69098 402 69119 458
rect 69175 402 69196 458
rect 69098 381 69196 402
rect 71594 458 71692 479
rect 71594 402 71615 458
rect 71671 402 71692 458
rect 71594 381 71692 402
rect 74090 458 74188 479
rect 74090 402 74111 458
rect 74167 402 74188 458
rect 74090 381 74188 402
rect 76586 458 76684 479
rect 76586 402 76607 458
rect 76663 402 76684 458
rect 76586 381 76684 402
rect 79082 458 79180 479
rect 79082 402 79103 458
rect 79159 402 79180 458
rect 79082 381 79180 402
rect 1706 136 1804 157
rect 1706 80 1727 136
rect 1783 80 1804 136
rect 1706 59 1804 80
rect 4202 136 4300 157
rect 4202 80 4223 136
rect 4279 80 4300 136
rect 4202 59 4300 80
rect 6698 136 6796 157
rect 6698 80 6719 136
rect 6775 80 6796 136
rect 6698 59 6796 80
rect 9194 136 9292 157
rect 9194 80 9215 136
rect 9271 80 9292 136
rect 9194 59 9292 80
rect 11690 136 11788 157
rect 11690 80 11711 136
rect 11767 80 11788 136
rect 11690 59 11788 80
rect 14186 136 14284 157
rect 14186 80 14207 136
rect 14263 80 14284 136
rect 14186 59 14284 80
rect 16682 136 16780 157
rect 16682 80 16703 136
rect 16759 80 16780 136
rect 16682 59 16780 80
rect 19178 136 19276 157
rect 19178 80 19199 136
rect 19255 80 19276 136
rect 19178 59 19276 80
rect 21674 136 21772 157
rect 21674 80 21695 136
rect 21751 80 21772 136
rect 21674 59 21772 80
rect 24170 136 24268 157
rect 24170 80 24191 136
rect 24247 80 24268 136
rect 24170 59 24268 80
rect 26666 136 26764 157
rect 26666 80 26687 136
rect 26743 80 26764 136
rect 26666 59 26764 80
rect 29162 136 29260 157
rect 29162 80 29183 136
rect 29239 80 29260 136
rect 29162 59 29260 80
rect 31658 136 31756 157
rect 31658 80 31679 136
rect 31735 80 31756 136
rect 31658 59 31756 80
rect 34154 136 34252 157
rect 34154 80 34175 136
rect 34231 80 34252 136
rect 34154 59 34252 80
rect 36650 136 36748 157
rect 36650 80 36671 136
rect 36727 80 36748 136
rect 36650 59 36748 80
rect 39146 136 39244 157
rect 39146 80 39167 136
rect 39223 80 39244 136
rect 39146 59 39244 80
rect 41642 136 41740 157
rect 41642 80 41663 136
rect 41719 80 41740 136
rect 41642 59 41740 80
rect 44138 136 44236 157
rect 44138 80 44159 136
rect 44215 80 44236 136
rect 44138 59 44236 80
rect 46634 136 46732 157
rect 46634 80 46655 136
rect 46711 80 46732 136
rect 46634 59 46732 80
rect 49130 136 49228 157
rect 49130 80 49151 136
rect 49207 80 49228 136
rect 49130 59 49228 80
rect 51626 136 51724 157
rect 51626 80 51647 136
rect 51703 80 51724 136
rect 51626 59 51724 80
rect 54122 136 54220 157
rect 54122 80 54143 136
rect 54199 80 54220 136
rect 54122 59 54220 80
rect 56618 136 56716 157
rect 56618 80 56639 136
rect 56695 80 56716 136
rect 56618 59 56716 80
rect 59114 136 59212 157
rect 59114 80 59135 136
rect 59191 80 59212 136
rect 59114 59 59212 80
rect 61610 136 61708 157
rect 61610 80 61631 136
rect 61687 80 61708 136
rect 61610 59 61708 80
rect 64106 136 64204 157
rect 64106 80 64127 136
rect 64183 80 64204 136
rect 64106 59 64204 80
rect 66602 136 66700 157
rect 66602 80 66623 136
rect 66679 80 66700 136
rect 66602 59 66700 80
rect 69098 136 69196 157
rect 69098 80 69119 136
rect 69175 80 69196 136
rect 69098 59 69196 80
rect 71594 136 71692 157
rect 71594 80 71615 136
rect 71671 80 71692 136
rect 71594 59 71692 80
rect 74090 136 74188 157
rect 74090 80 74111 136
rect 74167 80 74188 136
rect 74090 59 74188 80
rect 76586 136 76684 157
rect 76586 80 76607 136
rect 76663 80 76684 136
rect 76586 59 76684 80
rect 79082 136 79180 157
rect 79082 80 79103 136
rect 79159 80 79180 136
rect 79082 59 79180 80
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_0
timestamp 1683767628
transform 1 0 18846 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_1
timestamp 1683767628
transform 1 0 16350 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_2
timestamp 1683767628
transform 1 0 13854 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_3
timestamp 1683767628
transform 1 0 11358 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_4
timestamp 1683767628
transform 1 0 8862 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_5
timestamp 1683767628
transform 1 0 6366 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_6
timestamp 1683767628
transform 1 0 3870 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_7
timestamp 1683767628
transform 1 0 1374 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_8
timestamp 1683767628
transform 1 0 38814 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_9
timestamp 1683767628
transform 1 0 36318 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_10
timestamp 1683767628
transform 1 0 33822 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_11
timestamp 1683767628
transform 1 0 31326 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_12
timestamp 1683767628
transform 1 0 28830 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_13
timestamp 1683767628
transform 1 0 26334 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_14
timestamp 1683767628
transform 1 0 23838 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_15
timestamp 1683767628
transform 1 0 21342 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_16
timestamp 1683767628
transform 1 0 58782 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_17
timestamp 1683767628
transform 1 0 56286 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_18
timestamp 1683767628
transform 1 0 53790 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_19
timestamp 1683767628
transform 1 0 51294 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_20
timestamp 1683767628
transform 1 0 48798 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_21
timestamp 1683767628
transform 1 0 46302 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_22
timestamp 1683767628
transform 1 0 43806 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_23
timestamp 1683767628
transform 1 0 41310 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_24
timestamp 1683767628
transform 1 0 78750 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_25
timestamp 1683767628
transform 1 0 76254 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_26
timestamp 1683767628
transform 1 0 73758 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_27
timestamp 1683767628
transform 1 0 71262 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_28
timestamp 1683767628
transform 1 0 68766 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_29
timestamp 1683767628
transform 1 0 66270 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_30
timestamp 1683767628
transform 1 0 63774 0 1 0
box -541 0 937 2256
use sky130_fd_bd_sram__openram_sense_amp_2  sky130_fd_bd_sram__openram_sense_amp_31
timestamp 1683767628
transform 1 0 61278 0 1 0
box -541 0 937 2256
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_0
timestamp 1683767628
transform 1 0 6714 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_1
timestamp 1683767628
transform 1 0 6702 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_2
timestamp 1683767628
transform 1 0 6714 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_3
timestamp 1683767628
transform 1 0 6784 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_4
timestamp 1683767628
transform 1 0 4218 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_5
timestamp 1683767628
transform 1 0 4206 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_6
timestamp 1683767628
transform 1 0 4218 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_7
timestamp 1683767628
transform 1 0 4288 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_8
timestamp 1683767628
transform 1 0 1722 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_9
timestamp 1683767628
transform 1 0 1710 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_10
timestamp 1683767628
transform 1 0 1722 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_11
timestamp 1683767628
transform 1 0 1792 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_12
timestamp 1683767628
transform 1 0 19194 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_13
timestamp 1683767628
transform 1 0 19182 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_14
timestamp 1683767628
transform 1 0 19194 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_15
timestamp 1683767628
transform 1 0 19264 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_16
timestamp 1683767628
transform 1 0 16698 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_17
timestamp 1683767628
transform 1 0 16686 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_18
timestamp 1683767628
transform 1 0 16698 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_19
timestamp 1683767628
transform 1 0 16768 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_20
timestamp 1683767628
transform 1 0 18936 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_21
timestamp 1683767628
transform 1 0 16440 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_22
timestamp 1683767628
transform 1 0 13944 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_23
timestamp 1683767628
transform 1 0 11448 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_24
timestamp 1683767628
transform 1 0 8952 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_25
timestamp 1683767628
transform 1 0 6456 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_26
timestamp 1683767628
transform 1 0 3960 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_27
timestamp 1683767628
transform 1 0 1464 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_28
timestamp 1683767628
transform 1 0 14202 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_29
timestamp 1683767628
transform 1 0 14190 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_30
timestamp 1683767628
transform 1 0 14202 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_31
timestamp 1683767628
transform 1 0 14272 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_32
timestamp 1683767628
transform 1 0 11706 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_33
timestamp 1683767628
transform 1 0 11694 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_34
timestamp 1683767628
transform 1 0 11706 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_35
timestamp 1683767628
transform 1 0 11776 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_36
timestamp 1683767628
transform 1 0 9210 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_37
timestamp 1683767628
transform 1 0 9198 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_38
timestamp 1683767628
transform 1 0 9210 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_39
timestamp 1683767628
transform 1 0 9280 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_40
timestamp 1683767628
transform 1 0 39162 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_41
timestamp 1683767628
transform 1 0 39150 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_42
timestamp 1683767628
transform 1 0 39162 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_43
timestamp 1683767628
transform 1 0 39232 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_44
timestamp 1683767628
transform 1 0 36666 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_45
timestamp 1683767628
transform 1 0 36654 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_46
timestamp 1683767628
transform 1 0 36666 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_47
timestamp 1683767628
transform 1 0 36736 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_48
timestamp 1683767628
transform 1 0 38904 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_49
timestamp 1683767628
transform 1 0 36408 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_50
timestamp 1683767628
transform 1 0 33912 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_51
timestamp 1683767628
transform 1 0 31416 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_52
timestamp 1683767628
transform 1 0 28920 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_53
timestamp 1683767628
transform 1 0 26424 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_54
timestamp 1683767628
transform 1 0 23928 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_55
timestamp 1683767628
transform 1 0 21432 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_56
timestamp 1683767628
transform 1 0 34170 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_57
timestamp 1683767628
transform 1 0 34158 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_58
timestamp 1683767628
transform 1 0 34170 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_59
timestamp 1683767628
transform 1 0 34240 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_60
timestamp 1683767628
transform 1 0 31674 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_61
timestamp 1683767628
transform 1 0 31662 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_62
timestamp 1683767628
transform 1 0 31674 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_63
timestamp 1683767628
transform 1 0 31744 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_64
timestamp 1683767628
transform 1 0 29178 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_65
timestamp 1683767628
transform 1 0 29166 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_66
timestamp 1683767628
transform 1 0 29178 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_67
timestamp 1683767628
transform 1 0 29248 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_68
timestamp 1683767628
transform 1 0 26682 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_69
timestamp 1683767628
transform 1 0 26670 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_70
timestamp 1683767628
transform 1 0 26682 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_71
timestamp 1683767628
transform 1 0 26752 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_72
timestamp 1683767628
transform 1 0 24186 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_73
timestamp 1683767628
transform 1 0 24174 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_74
timestamp 1683767628
transform 1 0 24186 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_75
timestamp 1683767628
transform 1 0 24256 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_76
timestamp 1683767628
transform 1 0 21690 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_77
timestamp 1683767628
transform 1 0 21678 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_78
timestamp 1683767628
transform 1 0 21690 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_79
timestamp 1683767628
transform 1 0 21760 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_80
timestamp 1683767628
transform 1 0 59130 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_81
timestamp 1683767628
transform 1 0 59118 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_82
timestamp 1683767628
transform 1 0 59130 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_83
timestamp 1683767628
transform 1 0 59200 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_84
timestamp 1683767628
transform 1 0 58872 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_85
timestamp 1683767628
transform 1 0 56376 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_86
timestamp 1683767628
transform 1 0 53880 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_87
timestamp 1683767628
transform 1 0 51384 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_88
timestamp 1683767628
transform 1 0 48888 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_89
timestamp 1683767628
transform 1 0 46392 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_90
timestamp 1683767628
transform 1 0 43896 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_91
timestamp 1683767628
transform 1 0 41400 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_92
timestamp 1683767628
transform 1 0 56634 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_93
timestamp 1683767628
transform 1 0 56622 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_94
timestamp 1683767628
transform 1 0 56634 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_95
timestamp 1683767628
transform 1 0 56704 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_96
timestamp 1683767628
transform 1 0 54138 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_97
timestamp 1683767628
transform 1 0 54126 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_98
timestamp 1683767628
transform 1 0 54138 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_99
timestamp 1683767628
transform 1 0 54208 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_100
timestamp 1683767628
transform 1 0 51642 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_101
timestamp 1683767628
transform 1 0 51630 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_102
timestamp 1683767628
transform 1 0 51642 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_103
timestamp 1683767628
transform 1 0 51712 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_104
timestamp 1683767628
transform 1 0 49146 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_105
timestamp 1683767628
transform 1 0 49134 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_106
timestamp 1683767628
transform 1 0 49146 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_107
timestamp 1683767628
transform 1 0 49216 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_108
timestamp 1683767628
transform 1 0 46650 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_109
timestamp 1683767628
transform 1 0 46638 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_110
timestamp 1683767628
transform 1 0 46650 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_111
timestamp 1683767628
transform 1 0 46720 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_112
timestamp 1683767628
transform 1 0 44154 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_113
timestamp 1683767628
transform 1 0 44142 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_114
timestamp 1683767628
transform 1 0 44154 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_115
timestamp 1683767628
transform 1 0 44224 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_116
timestamp 1683767628
transform 1 0 41658 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_117
timestamp 1683767628
transform 1 0 41646 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_118
timestamp 1683767628
transform 1 0 41658 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_119
timestamp 1683767628
transform 1 0 41728 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_120
timestamp 1683767628
transform 1 0 78840 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_121
timestamp 1683767628
transform 1 0 76344 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_122
timestamp 1683767628
transform 1 0 73848 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_123
timestamp 1683767628
transform 1 0 71352 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_124
timestamp 1683767628
transform 1 0 68856 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_125
timestamp 1683767628
transform 1 0 66360 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_126
timestamp 1683767628
transform 1 0 63864 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_127
timestamp 1683767628
transform 1 0 61368 0 1 2157
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_128
timestamp 1683767628
transform 1 0 79098 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_129
timestamp 1683767628
transform 1 0 79086 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_130
timestamp 1683767628
transform 1 0 79098 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_131
timestamp 1683767628
transform 1 0 79168 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_132
timestamp 1683767628
transform 1 0 76602 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_133
timestamp 1683767628
transform 1 0 76590 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_134
timestamp 1683767628
transform 1 0 76602 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_135
timestamp 1683767628
transform 1 0 76672 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_136
timestamp 1683767628
transform 1 0 74106 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_137
timestamp 1683767628
transform 1 0 74094 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_138
timestamp 1683767628
transform 1 0 74106 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_139
timestamp 1683767628
transform 1 0 74176 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_140
timestamp 1683767628
transform 1 0 71610 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_141
timestamp 1683767628
transform 1 0 71598 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_142
timestamp 1683767628
transform 1 0 71610 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_143
timestamp 1683767628
transform 1 0 71680 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_144
timestamp 1683767628
transform 1 0 69114 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_145
timestamp 1683767628
transform 1 0 69102 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_146
timestamp 1683767628
transform 1 0 69114 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_147
timestamp 1683767628
transform 1 0 69184 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_148
timestamp 1683767628
transform 1 0 66618 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_149
timestamp 1683767628
transform 1 0 66606 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_150
timestamp 1683767628
transform 1 0 66618 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_151
timestamp 1683767628
transform 1 0 66688 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_152
timestamp 1683767628
transform 1 0 64122 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_153
timestamp 1683767628
transform 1 0 64110 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_154
timestamp 1683767628
transform 1 0 64122 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_155
timestamp 1683767628
transform 1 0 64192 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_156
timestamp 1683767628
transform 1 0 61626 0 1 393
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_157
timestamp 1683767628
transform 1 0 61614 0 1 1231
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_158
timestamp 1683767628
transform 1 0 61626 0 1 71
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_159
timestamp 1683767628
transform 1 0 61696 0 1 2005
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_0
timestamp 1683767628
transform 1 0 6715 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_1
timestamp 1683767628
transform 1 0 6703 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_2
timestamp 1683767628
transform 1 0 6715 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_3
timestamp 1683767628
transform 1 0 6785 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_4
timestamp 1683767628
transform 1 0 4219 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_5
timestamp 1683767628
transform 1 0 4207 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_6
timestamp 1683767628
transform 1 0 4219 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_7
timestamp 1683767628
transform 1 0 4289 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_8
timestamp 1683767628
transform 1 0 1723 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_9
timestamp 1683767628
transform 1 0 1711 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_10
timestamp 1683767628
transform 1 0 1723 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_11
timestamp 1683767628
transform 1 0 1793 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_12
timestamp 1683767628
transform 1 0 19195 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_13
timestamp 1683767628
transform 1 0 19183 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_14
timestamp 1683767628
transform 1 0 19195 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_15
timestamp 1683767628
transform 1 0 19265 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_16
timestamp 1683767628
transform 1 0 16699 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_17
timestamp 1683767628
transform 1 0 16687 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_18
timestamp 1683767628
transform 1 0 16699 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_19
timestamp 1683767628
transform 1 0 16769 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_20
timestamp 1683767628
transform 1 0 18937 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_21
timestamp 1683767628
transform 1 0 16441 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_22
timestamp 1683767628
transform 1 0 13945 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_23
timestamp 1683767628
transform 1 0 11449 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_24
timestamp 1683767628
transform 1 0 8953 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_25
timestamp 1683767628
transform 1 0 6457 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_26
timestamp 1683767628
transform 1 0 3961 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_27
timestamp 1683767628
transform 1 0 1465 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_28
timestamp 1683767628
transform 1 0 14203 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_29
timestamp 1683767628
transform 1 0 14191 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_30
timestamp 1683767628
transform 1 0 14203 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_31
timestamp 1683767628
transform 1 0 14273 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_32
timestamp 1683767628
transform 1 0 11707 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_33
timestamp 1683767628
transform 1 0 11695 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_34
timestamp 1683767628
transform 1 0 11707 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_35
timestamp 1683767628
transform 1 0 11777 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_36
timestamp 1683767628
transform 1 0 9211 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_37
timestamp 1683767628
transform 1 0 9199 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_38
timestamp 1683767628
transform 1 0 9211 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_39
timestamp 1683767628
transform 1 0 9281 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_40
timestamp 1683767628
transform 1 0 39163 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_41
timestamp 1683767628
transform 1 0 39151 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_42
timestamp 1683767628
transform 1 0 39163 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_43
timestamp 1683767628
transform 1 0 39233 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_44
timestamp 1683767628
transform 1 0 36667 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_45
timestamp 1683767628
transform 1 0 36655 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_46
timestamp 1683767628
transform 1 0 36667 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_47
timestamp 1683767628
transform 1 0 36737 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_48
timestamp 1683767628
transform 1 0 38905 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_49
timestamp 1683767628
transform 1 0 36409 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_50
timestamp 1683767628
transform 1 0 33913 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_51
timestamp 1683767628
transform 1 0 31417 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_52
timestamp 1683767628
transform 1 0 28921 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_53
timestamp 1683767628
transform 1 0 26425 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_54
timestamp 1683767628
transform 1 0 23929 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_55
timestamp 1683767628
transform 1 0 21433 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_56
timestamp 1683767628
transform 1 0 34171 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_57
timestamp 1683767628
transform 1 0 34159 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_58
timestamp 1683767628
transform 1 0 34171 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_59
timestamp 1683767628
transform 1 0 34241 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_60
timestamp 1683767628
transform 1 0 31675 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_61
timestamp 1683767628
transform 1 0 31663 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_62
timestamp 1683767628
transform 1 0 31675 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_63
timestamp 1683767628
transform 1 0 31745 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_64
timestamp 1683767628
transform 1 0 29179 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_65
timestamp 1683767628
transform 1 0 29167 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_66
timestamp 1683767628
transform 1 0 29179 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_67
timestamp 1683767628
transform 1 0 29249 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_68
timestamp 1683767628
transform 1 0 26683 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_69
timestamp 1683767628
transform 1 0 26671 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_70
timestamp 1683767628
transform 1 0 26683 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_71
timestamp 1683767628
transform 1 0 26753 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_72
timestamp 1683767628
transform 1 0 24187 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_73
timestamp 1683767628
transform 1 0 24175 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_74
timestamp 1683767628
transform 1 0 24187 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_75
timestamp 1683767628
transform 1 0 24257 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_76
timestamp 1683767628
transform 1 0 21691 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_77
timestamp 1683767628
transform 1 0 21679 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_78
timestamp 1683767628
transform 1 0 21691 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_79
timestamp 1683767628
transform 1 0 21761 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_80
timestamp 1683767628
transform 1 0 59131 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_81
timestamp 1683767628
transform 1 0 59119 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_82
timestamp 1683767628
transform 1 0 59131 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_83
timestamp 1683767628
transform 1 0 59201 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_84
timestamp 1683767628
transform 1 0 58873 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_85
timestamp 1683767628
transform 1 0 56377 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_86
timestamp 1683767628
transform 1 0 53881 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_87
timestamp 1683767628
transform 1 0 51385 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_88
timestamp 1683767628
transform 1 0 48889 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_89
timestamp 1683767628
transform 1 0 46393 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_90
timestamp 1683767628
transform 1 0 43897 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_91
timestamp 1683767628
transform 1 0 41401 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_92
timestamp 1683767628
transform 1 0 56635 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_93
timestamp 1683767628
transform 1 0 56623 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_94
timestamp 1683767628
transform 1 0 56635 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_95
timestamp 1683767628
transform 1 0 56705 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_96
timestamp 1683767628
transform 1 0 54139 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_97
timestamp 1683767628
transform 1 0 54127 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_98
timestamp 1683767628
transform 1 0 54139 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_99
timestamp 1683767628
transform 1 0 54209 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_100
timestamp 1683767628
transform 1 0 51643 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_101
timestamp 1683767628
transform 1 0 51631 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_102
timestamp 1683767628
transform 1 0 51643 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_103
timestamp 1683767628
transform 1 0 51713 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_104
timestamp 1683767628
transform 1 0 49147 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_105
timestamp 1683767628
transform 1 0 49135 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_106
timestamp 1683767628
transform 1 0 49147 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_107
timestamp 1683767628
transform 1 0 49217 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_108
timestamp 1683767628
transform 1 0 46651 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_109
timestamp 1683767628
transform 1 0 46639 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_110
timestamp 1683767628
transform 1 0 46651 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_111
timestamp 1683767628
transform 1 0 46721 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_112
timestamp 1683767628
transform 1 0 44155 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_113
timestamp 1683767628
transform 1 0 44143 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_114
timestamp 1683767628
transform 1 0 44155 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_115
timestamp 1683767628
transform 1 0 44225 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_116
timestamp 1683767628
transform 1 0 41659 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_117
timestamp 1683767628
transform 1 0 41647 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_118
timestamp 1683767628
transform 1 0 41659 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_119
timestamp 1683767628
transform 1 0 41729 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_120
timestamp 1683767628
transform 1 0 78841 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_121
timestamp 1683767628
transform 1 0 76345 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_122
timestamp 1683767628
transform 1 0 73849 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_123
timestamp 1683767628
transform 1 0 71353 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_124
timestamp 1683767628
transform 1 0 68857 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_125
timestamp 1683767628
transform 1 0 66361 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_126
timestamp 1683767628
transform 1 0 63865 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_127
timestamp 1683767628
transform 1 0 61369 0 1 2162
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_128
timestamp 1683767628
transform 1 0 79099 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_129
timestamp 1683767628
transform 1 0 79087 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_130
timestamp 1683767628
transform 1 0 79099 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_131
timestamp 1683767628
transform 1 0 79169 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_132
timestamp 1683767628
transform 1 0 76603 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_133
timestamp 1683767628
transform 1 0 76591 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_134
timestamp 1683767628
transform 1 0 76603 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_135
timestamp 1683767628
transform 1 0 76673 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_136
timestamp 1683767628
transform 1 0 74107 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_137
timestamp 1683767628
transform 1 0 74095 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_138
timestamp 1683767628
transform 1 0 74107 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_139
timestamp 1683767628
transform 1 0 74177 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_140
timestamp 1683767628
transform 1 0 71611 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_141
timestamp 1683767628
transform 1 0 71599 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_142
timestamp 1683767628
transform 1 0 71611 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_143
timestamp 1683767628
transform 1 0 71681 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_144
timestamp 1683767628
transform 1 0 69115 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_145
timestamp 1683767628
transform 1 0 69103 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_146
timestamp 1683767628
transform 1 0 69115 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_147
timestamp 1683767628
transform 1 0 69185 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_148
timestamp 1683767628
transform 1 0 66619 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_149
timestamp 1683767628
transform 1 0 66607 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_150
timestamp 1683767628
transform 1 0 66619 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_151
timestamp 1683767628
transform 1 0 66689 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_152
timestamp 1683767628
transform 1 0 64123 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_153
timestamp 1683767628
transform 1 0 64111 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_154
timestamp 1683767628
transform 1 0 64123 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_155
timestamp 1683767628
transform 1 0 64193 0 1 2010
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_156
timestamp 1683767628
transform 1 0 61627 0 1 398
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_157
timestamp 1683767628
transform 1 0 61615 0 1 1236
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_158
timestamp 1683767628
transform 1 0 61627 0 1 76
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_159
timestamp 1683767628
transform 1 0 61697 0 1 2010
box 0 0 1 1
<< labels >>
rlabel metal3 s 46704 1993 46802 2091 4 gnd
port 1 nsew
rlabel metal3 s 76656 1993 76754 2091 4 gnd
port 1 nsew
rlabel metal3 s 41712 1993 41810 2091 4 gnd
port 1 nsew
rlabel metal3 s 71664 1993 71762 2091 4 gnd
port 1 nsew
rlabel metal3 s 79152 1993 79250 2091 4 gnd
port 1 nsew
rlabel metal3 s 51696 1993 51794 2091 4 gnd
port 1 nsew
rlabel metal3 s 44208 1993 44306 2091 4 gnd
port 1 nsew
rlabel metal3 s 69168 1993 69266 2091 4 gnd
port 1 nsew
rlabel metal3 s 64176 1993 64274 2091 4 gnd
port 1 nsew
rlabel metal3 s 61680 1993 61778 2091 4 gnd
port 1 nsew
rlabel metal3 s 59184 1993 59282 2091 4 gnd
port 1 nsew
rlabel metal3 s 56688 1993 56786 2091 4 gnd
port 1 nsew
rlabel metal3 s 49200 1993 49298 2091 4 gnd
port 1 nsew
rlabel metal3 s 74160 1993 74258 2091 4 gnd
port 1 nsew
rlabel metal3 s 66672 1993 66770 2091 4 gnd
port 1 nsew
rlabel metal3 s 54192 1993 54290 2091 4 gnd
port 1 nsew
rlabel metal3 s 56618 381 56716 479 4 vdd
port 2 nsew
rlabel metal3 s 69086 1219 69184 1317 4 vdd
port 2 nsew
rlabel metal3 s 54122 381 54220 479 4 vdd
port 2 nsew
rlabel metal3 s 69098 381 69196 479 4 vdd
port 2 nsew
rlabel metal3 s 59102 1219 59200 1317 4 vdd
port 2 nsew
rlabel metal3 s 51614 1219 51712 1317 4 vdd
port 2 nsew
rlabel metal3 s 46634 381 46732 479 4 vdd
port 2 nsew
rlabel metal3 s 61610 381 61708 479 4 vdd
port 2 nsew
rlabel metal3 s 71582 1219 71680 1317 4 vdd
port 2 nsew
rlabel metal3 s 49130 381 49228 479 4 vdd
port 2 nsew
rlabel metal3 s 76586 381 76684 479 4 vdd
port 2 nsew
rlabel metal3 s 61598 1219 61696 1317 4 vdd
port 2 nsew
rlabel metal3 s 56606 1219 56704 1317 4 vdd
port 2 nsew
rlabel metal3 s 44138 381 44236 479 4 vdd
port 2 nsew
rlabel metal3 s 79070 1219 79168 1317 4 vdd
port 2 nsew
rlabel metal3 s 49118 1219 49216 1317 4 vdd
port 2 nsew
rlabel metal3 s 64106 381 64204 479 4 vdd
port 2 nsew
rlabel metal3 s 41630 1219 41728 1317 4 vdd
port 2 nsew
rlabel metal3 s 71594 381 71692 479 4 vdd
port 2 nsew
rlabel metal3 s 54110 1219 54208 1317 4 vdd
port 2 nsew
rlabel metal3 s 44126 1219 44224 1317 4 vdd
port 2 nsew
rlabel metal3 s 76574 1219 76672 1317 4 vdd
port 2 nsew
rlabel metal3 s 74078 1219 74176 1317 4 vdd
port 2 nsew
rlabel metal3 s 74090 381 74188 479 4 vdd
port 2 nsew
rlabel metal3 s 66602 381 66700 479 4 vdd
port 2 nsew
rlabel metal3 s 59114 381 59212 479 4 vdd
port 2 nsew
rlabel metal3 s 41642 381 41740 479 4 vdd
port 2 nsew
rlabel metal3 s 46622 1219 46720 1317 4 vdd
port 2 nsew
rlabel metal3 s 64094 1219 64192 1317 4 vdd
port 2 nsew
rlabel metal3 s 66590 1219 66688 1317 4 vdd
port 2 nsew
rlabel metal3 s 79082 381 79180 479 4 vdd
port 2 nsew
rlabel metal3 s 51626 381 51724 479 4 vdd
port 2 nsew
rlabel metal3 s 9264 1993 9362 2091 4 gnd
port 1 nsew
rlabel metal3 s 14186 381 14284 479 4 vdd
port 2 nsew
rlabel metal3 s 21744 1993 21842 2091 4 gnd
port 1 nsew
rlabel metal3 s 34224 1993 34322 2091 4 gnd
port 1 nsew
rlabel metal3 s 39216 1993 39314 2091 4 gnd
port 1 nsew
rlabel metal3 s 16752 1993 16850 2091 4 gnd
port 1 nsew
rlabel metal3 s 4272 1993 4370 2091 4 gnd
port 1 nsew
rlabel metal3 s 36650 381 36748 479 4 vdd
port 2 nsew
rlabel metal3 s 11760 1993 11858 2091 4 gnd
port 1 nsew
rlabel metal3 s 36720 1993 36818 2091 4 gnd
port 1 nsew
rlabel metal3 s 24240 1993 24338 2091 4 gnd
port 1 nsew
rlabel metal3 s 31658 381 31756 479 4 vdd
port 2 nsew
rlabel metal3 s 14174 1219 14272 1317 4 vdd
port 2 nsew
rlabel metal3 s 29232 1993 29330 2091 4 gnd
port 1 nsew
rlabel metal3 s 26654 1219 26752 1317 4 vdd
port 2 nsew
rlabel metal3 s 14256 1993 14354 2091 4 gnd
port 1 nsew
rlabel metal3 s 36638 1219 36736 1317 4 vdd
port 2 nsew
rlabel metal3 s 16682 381 16780 479 4 vdd
port 2 nsew
rlabel metal3 s 1694 1219 1792 1317 4 vdd
port 2 nsew
rlabel metal3 s 1776 1993 1874 2091 4 gnd
port 1 nsew
rlabel metal3 s 21662 1219 21760 1317 4 vdd
port 2 nsew
rlabel metal3 s 31728 1993 31826 2091 4 gnd
port 1 nsew
rlabel metal3 s 24158 1219 24256 1317 4 vdd
port 2 nsew
rlabel metal3 s 31646 1219 31744 1317 4 vdd
port 2 nsew
rlabel metal3 s 4202 381 4300 479 4 vdd
port 2 nsew
rlabel metal3 s 39134 1219 39232 1317 4 vdd
port 2 nsew
rlabel metal3 s 11678 1219 11776 1317 4 vdd
port 2 nsew
rlabel metal3 s 34142 1219 34240 1317 4 vdd
port 2 nsew
rlabel metal3 s 29162 381 29260 479 4 vdd
port 2 nsew
rlabel metal3 s 19178 381 19276 479 4 vdd
port 2 nsew
rlabel metal3 s 19166 1219 19264 1317 4 vdd
port 2 nsew
rlabel metal3 s 6686 1219 6784 1317 4 vdd
port 2 nsew
rlabel metal3 s 24170 381 24268 479 4 vdd
port 2 nsew
rlabel metal3 s 39146 381 39244 479 4 vdd
port 2 nsew
rlabel metal3 s 11690 381 11788 479 4 vdd
port 2 nsew
rlabel metal3 s 4190 1219 4288 1317 4 vdd
port 2 nsew
rlabel metal3 s 9182 1219 9280 1317 4 vdd
port 2 nsew
rlabel metal3 s 6698 381 6796 479 4 vdd
port 2 nsew
rlabel metal3 s 21674 381 21772 479 4 vdd
port 2 nsew
rlabel metal3 s 34154 381 34252 479 4 vdd
port 2 nsew
rlabel metal3 s 1706 381 1804 479 4 vdd
port 2 nsew
rlabel metal3 s 26736 1993 26834 2091 4 gnd
port 1 nsew
rlabel metal3 s 19248 1993 19346 2091 4 gnd
port 1 nsew
rlabel metal3 s 26666 381 26764 479 4 vdd
port 2 nsew
rlabel metal3 s 6768 1993 6866 2091 4 gnd
port 1 nsew
rlabel metal3 s 9194 381 9292 479 4 vdd
port 2 nsew
rlabel metal3 s 16670 1219 16768 1317 4 vdd
port 2 nsew
rlabel metal3 s 29150 1219 29248 1317 4 vdd
port 2 nsew
rlabel metal3 s 0 2164 79250 2224 4 en
port 3 nsew
rlabel metal3 s 4202 59 4300 157 4 gnd
port 1 nsew
rlabel metal3 s 1706 59 1804 157 4 gnd
port 1 nsew
rlabel metal3 s 34154 59 34252 157 4 gnd
port 1 nsew
rlabel metal3 s 29162 59 29260 157 4 gnd
port 1 nsew
rlabel metal3 s 19178 59 19276 157 4 gnd
port 1 nsew
rlabel metal3 s 36650 59 36748 157 4 gnd
port 1 nsew
rlabel metal3 s 16682 59 16780 157 4 gnd
port 1 nsew
rlabel metal3 s 39146 59 39244 157 4 gnd
port 1 nsew
rlabel metal3 s 24170 59 24268 157 4 gnd
port 1 nsew
rlabel metal3 s 6698 59 6796 157 4 gnd
port 1 nsew
rlabel metal3 s 9194 59 9292 157 4 gnd
port 1 nsew
rlabel metal3 s 26666 59 26764 157 4 gnd
port 1 nsew
rlabel metal3 s 14186 59 14284 157 4 gnd
port 1 nsew
rlabel metal3 s 21674 59 21772 157 4 gnd
port 1 nsew
rlabel metal3 s 11690 59 11788 157 4 gnd
port 1 nsew
rlabel metal3 s 31658 59 31756 157 4 gnd
port 1 nsew
rlabel metal3 s 44138 59 44236 157 4 gnd
port 1 nsew
rlabel metal3 s 79082 59 79180 157 4 gnd
port 1 nsew
rlabel metal3 s 61610 59 61708 157 4 gnd
port 1 nsew
rlabel metal3 s 76586 59 76684 157 4 gnd
port 1 nsew
rlabel metal3 s 64106 59 64204 157 4 gnd
port 1 nsew
rlabel metal3 s 69098 59 69196 157 4 gnd
port 1 nsew
rlabel metal3 s 59114 59 59212 157 4 gnd
port 1 nsew
rlabel metal3 s 54122 59 54220 157 4 gnd
port 1 nsew
rlabel metal3 s 41642 59 41740 157 4 gnd
port 1 nsew
rlabel metal3 s 46634 59 46732 157 4 gnd
port 1 nsew
rlabel metal3 s 71594 59 71692 157 4 gnd
port 1 nsew
rlabel metal3 s 66602 59 66700 157 4 gnd
port 1 nsew
rlabel metal3 s 74090 59 74188 157 4 gnd
port 1 nsew
rlabel metal3 s 49130 59 49228 157 4 gnd
port 1 nsew
rlabel metal3 s 51626 59 51724 157 4 gnd
port 1 nsew
rlabel metal3 s 56618 59 56716 157 4 gnd
port 1 nsew
rlabel metal1 s 1570 1130 1604 2256 4 bl_0
port 4 nsew
rlabel metal1 s 1646 1142 1674 2256 4 br_0
port 5 nsew
rlabel metal1 s 1478 0 1524 254 4 data_0
port 6 nsew
rlabel metal1 s 4066 1130 4100 2256 4 bl_1
port 7 nsew
rlabel metal1 s 4142 1142 4170 2256 4 br_1
port 8 nsew
rlabel metal1 s 3974 0 4020 254 4 data_1
port 9 nsew
rlabel metal1 s 6562 1130 6596 2256 4 bl_2
port 10 nsew
rlabel metal1 s 6638 1142 6666 2256 4 br_2
port 11 nsew
rlabel metal1 s 6470 0 6516 254 4 data_2
port 12 nsew
rlabel metal1 s 9058 1130 9092 2256 4 bl_3
port 13 nsew
rlabel metal1 s 9134 1142 9162 2256 4 br_3
port 14 nsew
rlabel metal1 s 8966 0 9012 254 4 data_3
port 15 nsew
rlabel metal1 s 11554 1130 11588 2256 4 bl_4
port 16 nsew
rlabel metal1 s 11630 1142 11658 2256 4 br_4
port 17 nsew
rlabel metal1 s 11462 0 11508 254 4 data_4
port 18 nsew
rlabel metal1 s 14050 1130 14084 2256 4 bl_5
port 19 nsew
rlabel metal1 s 14126 1142 14154 2256 4 br_5
port 20 nsew
rlabel metal1 s 13958 0 14004 254 4 data_5
port 21 nsew
rlabel metal1 s 16546 1130 16580 2256 4 bl_6
port 22 nsew
rlabel metal1 s 16622 1142 16650 2256 4 br_6
port 23 nsew
rlabel metal1 s 16454 0 16500 254 4 data_6
port 24 nsew
rlabel metal1 s 19042 1130 19076 2256 4 bl_7
port 25 nsew
rlabel metal1 s 19118 1142 19146 2256 4 br_7
port 26 nsew
rlabel metal1 s 18950 0 18996 254 4 data_7
port 27 nsew
rlabel metal1 s 21538 1130 21572 2256 4 bl_8
port 28 nsew
rlabel metal1 s 21614 1142 21642 2256 4 br_8
port 29 nsew
rlabel metal1 s 21446 0 21492 254 4 data_8
port 30 nsew
rlabel metal1 s 24034 1130 24068 2256 4 bl_9
port 31 nsew
rlabel metal1 s 24110 1142 24138 2256 4 br_9
port 32 nsew
rlabel metal1 s 23942 0 23988 254 4 data_9
port 33 nsew
rlabel metal1 s 26530 1130 26564 2256 4 bl_10
port 34 nsew
rlabel metal1 s 26606 1142 26634 2256 4 br_10
port 35 nsew
rlabel metal1 s 26438 0 26484 254 4 data_10
port 36 nsew
rlabel metal1 s 29026 1130 29060 2256 4 bl_11
port 37 nsew
rlabel metal1 s 29102 1142 29130 2256 4 br_11
port 38 nsew
rlabel metal1 s 28934 0 28980 254 4 data_11
port 39 nsew
rlabel metal1 s 31522 1130 31556 2256 4 bl_12
port 40 nsew
rlabel metal1 s 31598 1142 31626 2256 4 br_12
port 41 nsew
rlabel metal1 s 31430 0 31476 254 4 data_12
port 42 nsew
rlabel metal1 s 34018 1130 34052 2256 4 bl_13
port 43 nsew
rlabel metal1 s 34094 1142 34122 2256 4 br_13
port 44 nsew
rlabel metal1 s 33926 0 33972 254 4 data_13
port 45 nsew
rlabel metal1 s 36514 1130 36548 2256 4 bl_14
port 46 nsew
rlabel metal1 s 36590 1142 36618 2256 4 br_14
port 47 nsew
rlabel metal1 s 36422 0 36468 254 4 data_14
port 48 nsew
rlabel metal1 s 39010 1130 39044 2256 4 bl_15
port 49 nsew
rlabel metal1 s 39086 1142 39114 2256 4 br_15
port 50 nsew
rlabel metal1 s 38918 0 38964 254 4 data_15
port 51 nsew
rlabel metal1 s 41506 1130 41540 2256 4 bl_16
port 52 nsew
rlabel metal1 s 41582 1142 41610 2256 4 br_16
port 53 nsew
rlabel metal1 s 41414 0 41460 254 4 data_16
port 54 nsew
rlabel metal1 s 44002 1130 44036 2256 4 bl_17
port 55 nsew
rlabel metal1 s 44078 1142 44106 2256 4 br_17
port 56 nsew
rlabel metal1 s 43910 0 43956 254 4 data_17
port 57 nsew
rlabel metal1 s 46498 1130 46532 2256 4 bl_18
port 58 nsew
rlabel metal1 s 46574 1142 46602 2256 4 br_18
port 59 nsew
rlabel metal1 s 46406 0 46452 254 4 data_18
port 60 nsew
rlabel metal1 s 48994 1130 49028 2256 4 bl_19
port 61 nsew
rlabel metal1 s 49070 1142 49098 2256 4 br_19
port 62 nsew
rlabel metal1 s 48902 0 48948 254 4 data_19
port 63 nsew
rlabel metal1 s 51490 1130 51524 2256 4 bl_20
port 64 nsew
rlabel metal1 s 51566 1142 51594 2256 4 br_20
port 65 nsew
rlabel metal1 s 51398 0 51444 254 4 data_20
port 66 nsew
rlabel metal1 s 53986 1130 54020 2256 4 bl_21
port 67 nsew
rlabel metal1 s 54062 1142 54090 2256 4 br_21
port 68 nsew
rlabel metal1 s 53894 0 53940 254 4 data_21
port 69 nsew
rlabel metal1 s 56482 1130 56516 2256 4 bl_22
port 70 nsew
rlabel metal1 s 56558 1142 56586 2256 4 br_22
port 71 nsew
rlabel metal1 s 56390 0 56436 254 4 data_22
port 72 nsew
rlabel metal1 s 58978 1130 59012 2256 4 bl_23
port 73 nsew
rlabel metal1 s 59054 1142 59082 2256 4 br_23
port 74 nsew
rlabel metal1 s 58886 0 58932 254 4 data_23
port 75 nsew
rlabel metal1 s 61474 1130 61508 2256 4 bl_24
port 76 nsew
rlabel metal1 s 61550 1142 61578 2256 4 br_24
port 77 nsew
rlabel metal1 s 61382 0 61428 254 4 data_24
port 78 nsew
rlabel metal1 s 63970 1130 64004 2256 4 bl_25
port 79 nsew
rlabel metal1 s 64046 1142 64074 2256 4 br_25
port 80 nsew
rlabel metal1 s 63878 0 63924 254 4 data_25
port 81 nsew
rlabel metal1 s 66466 1130 66500 2256 4 bl_26
port 82 nsew
rlabel metal1 s 66542 1142 66570 2256 4 br_26
port 83 nsew
rlabel metal1 s 66374 0 66420 254 4 data_26
port 84 nsew
rlabel metal1 s 68962 1130 68996 2256 4 bl_27
port 85 nsew
rlabel metal1 s 69038 1142 69066 2256 4 br_27
port 86 nsew
rlabel metal1 s 68870 0 68916 254 4 data_27
port 87 nsew
rlabel metal1 s 71458 1130 71492 2256 4 bl_28
port 88 nsew
rlabel metal1 s 71534 1142 71562 2256 4 br_28
port 89 nsew
rlabel metal1 s 71366 0 71412 254 4 data_28
port 90 nsew
rlabel metal1 s 73954 1130 73988 2256 4 bl_29
port 91 nsew
rlabel metal1 s 74030 1142 74058 2256 4 br_29
port 92 nsew
rlabel metal1 s 73862 0 73908 254 4 data_29
port 93 nsew
rlabel metal1 s 76450 1130 76484 2256 4 bl_30
port 94 nsew
rlabel metal1 s 76526 1142 76554 2256 4 br_30
port 95 nsew
rlabel metal1 s 76358 0 76404 254 4 data_30
port 96 nsew
rlabel metal1 s 78946 1130 78980 2256 4 bl_31
port 97 nsew
rlabel metal1 s 79022 1142 79050 2256 4 br_31
port 98 nsew
rlabel metal1 s 78854 0 78900 254 4 data_31
port 99 nsew
<< properties >>
string FIXED_BBOX 0 0 79250 2256
string GDS_END 1522026
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 1446518
<< end >>
