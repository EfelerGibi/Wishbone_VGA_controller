magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect 576 2563 1795 3645
rect 576 2440 1648 2563
rect 576 1462 1817 2076
<< pwell >>
rect 186 569 2562 821
rect 204 415 2562 569
rect 1270 99 2562 415
rect 176 -231 2562 99
rect 176 -255 2522 -231
rect 146 -341 2522 -255
<< nmos >>
rect 255 -127 305 73
rect 361 -127 411 73
rect 467 -127 517 73
rect 683 -127 733 73
rect 789 -127 839 73
rect 895 -127 945 73
rect 1001 -127 1051 73
rect 1107 -127 1157 73
<< pmos >>
rect 1412 3491 1612 3541
rect 612 3385 1212 3435
rect 1412 3385 1612 3435
rect 612 3169 1612 3219
rect 612 3063 1612 3113
rect 612 2847 1612 2897
rect 612 2741 1612 2791
rect 612 2635 1612 2685
rect 612 2529 1612 2579
<< mvnmos >>
rect 265 595 425 795
rect 591 595 751 795
rect 807 595 967 795
rect 1023 595 1183 795
rect 1349 -205 1509 795
rect 1565 -205 1725 795
rect 1781 -205 1941 795
rect 1997 -205 2157 795
rect 2323 -205 2483 795
<< mvpmos >>
rect 642 1797 1642 1957
rect 642 1581 1642 1741
<< ndiff >>
rect 202 61 255 73
rect 202 27 210 61
rect 244 27 255 61
rect 202 -7 255 27
rect 202 -41 210 -7
rect 244 -41 255 -7
rect 202 -75 255 -41
rect 202 -109 210 -75
rect 244 -109 255 -75
rect 202 -127 255 -109
rect 305 61 361 73
rect 305 27 316 61
rect 350 27 361 61
rect 305 -7 361 27
rect 305 -41 316 -7
rect 350 -41 361 -7
rect 305 -75 361 -41
rect 305 -109 316 -75
rect 350 -109 361 -75
rect 305 -127 361 -109
rect 411 61 467 73
rect 411 27 422 61
rect 456 27 467 61
rect 411 -7 467 27
rect 411 -41 422 -7
rect 456 -41 467 -7
rect 411 -75 467 -41
rect 411 -109 422 -75
rect 456 -109 467 -75
rect 411 -127 467 -109
rect 517 61 570 73
rect 517 27 528 61
rect 562 27 570 61
rect 517 -7 570 27
rect 517 -41 528 -7
rect 562 -41 570 -7
rect 517 -75 570 -41
rect 517 -109 528 -75
rect 562 -109 570 -75
rect 517 -127 570 -109
rect 630 61 683 73
rect 630 27 638 61
rect 672 27 683 61
rect 630 -7 683 27
rect 630 -41 638 -7
rect 672 -41 683 -7
rect 630 -75 683 -41
rect 630 -109 638 -75
rect 672 -109 683 -75
rect 630 -127 683 -109
rect 733 61 789 73
rect 733 27 744 61
rect 778 27 789 61
rect 733 -7 789 27
rect 733 -41 744 -7
rect 778 -41 789 -7
rect 733 -75 789 -41
rect 733 -109 744 -75
rect 778 -109 789 -75
rect 733 -127 789 -109
rect 839 61 895 73
rect 839 27 850 61
rect 884 27 895 61
rect 839 -7 895 27
rect 839 -41 850 -7
rect 884 -41 895 -7
rect 839 -75 895 -41
rect 839 -109 850 -75
rect 884 -109 895 -75
rect 839 -127 895 -109
rect 945 61 1001 73
rect 945 27 956 61
rect 990 27 1001 61
rect 945 -7 1001 27
rect 945 -41 956 -7
rect 990 -41 1001 -7
rect 945 -75 1001 -41
rect 945 -109 956 -75
rect 990 -109 1001 -75
rect 945 -127 1001 -109
rect 1051 61 1107 73
rect 1051 27 1062 61
rect 1096 27 1107 61
rect 1051 -7 1107 27
rect 1051 -41 1062 -7
rect 1096 -41 1107 -7
rect 1051 -75 1107 -41
rect 1051 -109 1062 -75
rect 1096 -109 1107 -75
rect 1051 -127 1107 -109
rect 1157 61 1210 73
rect 1157 27 1168 61
rect 1202 27 1210 61
rect 1157 -7 1210 27
rect 1157 -41 1168 -7
rect 1202 -41 1210 -7
rect 1157 -75 1210 -41
rect 1157 -109 1168 -75
rect 1202 -109 1210 -75
rect 1157 -127 1210 -109
<< pdiff >>
rect 1412 3586 1612 3594
rect 1412 3552 1430 3586
rect 1464 3552 1498 3586
rect 1532 3552 1566 3586
rect 1600 3552 1612 3586
rect 1412 3541 1612 3552
rect 612 3480 1212 3488
rect 612 3446 690 3480
rect 724 3446 758 3480
rect 792 3446 826 3480
rect 860 3446 894 3480
rect 928 3446 962 3480
rect 996 3446 1030 3480
rect 1064 3446 1098 3480
rect 1132 3446 1166 3480
rect 1200 3446 1212 3480
rect 612 3435 1212 3446
rect 1412 3480 1612 3491
rect 1412 3446 1430 3480
rect 1464 3446 1498 3480
rect 1532 3446 1566 3480
rect 1600 3446 1612 3480
rect 1412 3435 1612 3446
rect 612 3374 1212 3385
rect 612 3340 690 3374
rect 724 3340 758 3374
rect 792 3340 826 3374
rect 860 3340 894 3374
rect 928 3340 962 3374
rect 996 3340 1030 3374
rect 1064 3340 1098 3374
rect 1132 3340 1166 3374
rect 1200 3340 1212 3374
rect 612 3332 1212 3340
rect 1412 3374 1612 3385
rect 1412 3340 1430 3374
rect 1464 3340 1498 3374
rect 1532 3340 1566 3374
rect 1600 3340 1612 3374
rect 1412 3332 1612 3340
rect 612 3264 1612 3272
rect 612 3230 682 3264
rect 716 3230 750 3264
rect 784 3230 818 3264
rect 852 3230 886 3264
rect 920 3230 954 3264
rect 988 3230 1022 3264
rect 1056 3230 1090 3264
rect 1124 3230 1158 3264
rect 1192 3230 1226 3264
rect 1260 3230 1294 3264
rect 1328 3230 1362 3264
rect 1396 3230 1430 3264
rect 1464 3230 1498 3264
rect 1532 3230 1566 3264
rect 1600 3230 1612 3264
rect 612 3219 1612 3230
rect 612 3158 1612 3169
rect 612 3124 682 3158
rect 716 3124 750 3158
rect 784 3124 818 3158
rect 852 3124 886 3158
rect 920 3124 954 3158
rect 988 3124 1022 3158
rect 1056 3124 1090 3158
rect 1124 3124 1158 3158
rect 1192 3124 1226 3158
rect 1260 3124 1294 3158
rect 1328 3124 1362 3158
rect 1396 3124 1430 3158
rect 1464 3124 1498 3158
rect 1532 3124 1566 3158
rect 1600 3124 1612 3158
rect 612 3113 1612 3124
rect 612 3052 1612 3063
rect 612 3018 682 3052
rect 716 3018 750 3052
rect 784 3018 818 3052
rect 852 3018 886 3052
rect 920 3018 954 3052
rect 988 3018 1022 3052
rect 1056 3018 1090 3052
rect 1124 3018 1158 3052
rect 1192 3018 1226 3052
rect 1260 3018 1294 3052
rect 1328 3018 1362 3052
rect 1396 3018 1430 3052
rect 1464 3018 1498 3052
rect 1532 3018 1566 3052
rect 1600 3018 1612 3052
rect 612 3010 1612 3018
rect 612 2942 1612 2950
rect 612 2908 682 2942
rect 716 2908 750 2942
rect 784 2908 818 2942
rect 852 2908 886 2942
rect 920 2908 954 2942
rect 988 2908 1022 2942
rect 1056 2908 1090 2942
rect 1124 2908 1158 2942
rect 1192 2908 1226 2942
rect 1260 2908 1294 2942
rect 1328 2908 1362 2942
rect 1396 2908 1430 2942
rect 1464 2908 1498 2942
rect 1532 2908 1566 2942
rect 1600 2908 1612 2942
rect 612 2897 1612 2908
rect 612 2836 1612 2847
rect 612 2802 682 2836
rect 716 2802 750 2836
rect 784 2802 818 2836
rect 852 2802 886 2836
rect 920 2802 954 2836
rect 988 2802 1022 2836
rect 1056 2802 1090 2836
rect 1124 2802 1158 2836
rect 1192 2802 1226 2836
rect 1260 2802 1294 2836
rect 1328 2802 1362 2836
rect 1396 2802 1430 2836
rect 1464 2802 1498 2836
rect 1532 2802 1566 2836
rect 1600 2802 1612 2836
rect 612 2791 1612 2802
rect 612 2730 1612 2741
rect 612 2696 682 2730
rect 716 2696 750 2730
rect 784 2696 818 2730
rect 852 2696 886 2730
rect 920 2696 954 2730
rect 988 2696 1022 2730
rect 1056 2696 1090 2730
rect 1124 2696 1158 2730
rect 1192 2696 1226 2730
rect 1260 2696 1294 2730
rect 1328 2696 1362 2730
rect 1396 2696 1430 2730
rect 1464 2696 1498 2730
rect 1532 2696 1566 2730
rect 1600 2696 1612 2730
rect 612 2685 1612 2696
rect 612 2624 1612 2635
rect 612 2590 682 2624
rect 716 2590 750 2624
rect 784 2590 818 2624
rect 852 2590 886 2624
rect 920 2590 954 2624
rect 988 2590 1022 2624
rect 1056 2590 1090 2624
rect 1124 2590 1158 2624
rect 1192 2590 1226 2624
rect 1260 2590 1294 2624
rect 1328 2590 1362 2624
rect 1396 2590 1430 2624
rect 1464 2590 1498 2624
rect 1532 2590 1566 2624
rect 1600 2590 1612 2624
rect 612 2579 1612 2590
rect 612 2518 1612 2529
rect 612 2484 682 2518
rect 716 2484 750 2518
rect 784 2484 818 2518
rect 852 2484 886 2518
rect 920 2484 954 2518
rect 988 2484 1022 2518
rect 1056 2484 1090 2518
rect 1124 2484 1158 2518
rect 1192 2484 1226 2518
rect 1260 2484 1294 2518
rect 1328 2484 1362 2518
rect 1396 2484 1430 2518
rect 1464 2484 1498 2518
rect 1532 2484 1566 2518
rect 1600 2484 1612 2518
rect 612 2476 1612 2484
<< mvndiff >>
rect 212 777 265 795
rect 212 743 220 777
rect 254 743 265 777
rect 212 709 265 743
rect 212 675 220 709
rect 254 675 265 709
rect 212 641 265 675
rect 212 607 220 641
rect 254 607 265 641
rect 212 595 265 607
rect 425 777 478 795
rect 425 743 436 777
rect 470 743 478 777
rect 425 709 478 743
rect 425 675 436 709
rect 470 675 478 709
rect 425 641 478 675
rect 425 607 436 641
rect 470 607 478 641
rect 425 595 478 607
rect 538 777 591 795
rect 538 743 546 777
rect 580 743 591 777
rect 538 709 591 743
rect 538 675 546 709
rect 580 675 591 709
rect 538 641 591 675
rect 538 607 546 641
rect 580 607 591 641
rect 538 595 591 607
rect 751 777 807 795
rect 751 743 762 777
rect 796 743 807 777
rect 751 709 807 743
rect 751 675 762 709
rect 796 675 807 709
rect 751 641 807 675
rect 751 607 762 641
rect 796 607 807 641
rect 751 595 807 607
rect 967 777 1023 795
rect 967 743 978 777
rect 1012 743 1023 777
rect 967 709 1023 743
rect 967 675 978 709
rect 1012 675 1023 709
rect 967 641 1023 675
rect 967 607 978 641
rect 1012 607 1023 641
rect 967 595 1023 607
rect 1183 777 1236 795
rect 1183 743 1194 777
rect 1228 743 1236 777
rect 1183 709 1236 743
rect 1183 675 1194 709
rect 1228 675 1236 709
rect 1183 641 1236 675
rect 1183 607 1194 641
rect 1228 607 1236 641
rect 1183 595 1236 607
rect 1296 725 1349 795
rect 1296 691 1304 725
rect 1338 691 1349 725
rect 1296 657 1349 691
rect 1296 623 1304 657
rect 1338 623 1349 657
rect 1296 589 1349 623
rect 1296 555 1304 589
rect 1338 555 1349 589
rect 1296 521 1349 555
rect 1296 487 1304 521
rect 1338 487 1349 521
rect 1296 453 1349 487
rect 1296 419 1304 453
rect 1338 419 1349 453
rect 1296 385 1349 419
rect 1296 351 1304 385
rect 1338 351 1349 385
rect 1296 317 1349 351
rect 1296 283 1304 317
rect 1338 283 1349 317
rect 1296 249 1349 283
rect 1296 215 1304 249
rect 1338 215 1349 249
rect 1296 181 1349 215
rect 1296 147 1304 181
rect 1338 147 1349 181
rect 1296 113 1349 147
rect 1296 79 1304 113
rect 1338 79 1349 113
rect 1296 45 1349 79
rect 1296 11 1304 45
rect 1338 11 1349 45
rect 1296 -23 1349 11
rect 1296 -57 1304 -23
rect 1338 -57 1349 -23
rect 1296 -91 1349 -57
rect 1296 -125 1304 -91
rect 1338 -125 1349 -91
rect 1296 -159 1349 -125
rect 1296 -193 1304 -159
rect 1338 -193 1349 -159
rect 1296 -205 1349 -193
rect 1509 725 1565 795
rect 1509 691 1520 725
rect 1554 691 1565 725
rect 1509 657 1565 691
rect 1509 623 1520 657
rect 1554 623 1565 657
rect 1509 589 1565 623
rect 1509 555 1520 589
rect 1554 555 1565 589
rect 1509 521 1565 555
rect 1509 487 1520 521
rect 1554 487 1565 521
rect 1509 453 1565 487
rect 1509 419 1520 453
rect 1554 419 1565 453
rect 1509 385 1565 419
rect 1509 351 1520 385
rect 1554 351 1565 385
rect 1509 317 1565 351
rect 1509 283 1520 317
rect 1554 283 1565 317
rect 1509 249 1565 283
rect 1509 215 1520 249
rect 1554 215 1565 249
rect 1509 181 1565 215
rect 1509 147 1520 181
rect 1554 147 1565 181
rect 1509 113 1565 147
rect 1509 79 1520 113
rect 1554 79 1565 113
rect 1509 45 1565 79
rect 1509 11 1520 45
rect 1554 11 1565 45
rect 1509 -23 1565 11
rect 1509 -57 1520 -23
rect 1554 -57 1565 -23
rect 1509 -91 1565 -57
rect 1509 -125 1520 -91
rect 1554 -125 1565 -91
rect 1509 -159 1565 -125
rect 1509 -193 1520 -159
rect 1554 -193 1565 -159
rect 1509 -205 1565 -193
rect 1725 725 1781 795
rect 1725 691 1736 725
rect 1770 691 1781 725
rect 1725 657 1781 691
rect 1725 623 1736 657
rect 1770 623 1781 657
rect 1725 589 1781 623
rect 1725 555 1736 589
rect 1770 555 1781 589
rect 1725 521 1781 555
rect 1725 487 1736 521
rect 1770 487 1781 521
rect 1725 453 1781 487
rect 1725 419 1736 453
rect 1770 419 1781 453
rect 1725 385 1781 419
rect 1725 351 1736 385
rect 1770 351 1781 385
rect 1725 317 1781 351
rect 1725 283 1736 317
rect 1770 283 1781 317
rect 1725 249 1781 283
rect 1725 215 1736 249
rect 1770 215 1781 249
rect 1725 181 1781 215
rect 1725 147 1736 181
rect 1770 147 1781 181
rect 1725 113 1781 147
rect 1725 79 1736 113
rect 1770 79 1781 113
rect 1725 45 1781 79
rect 1725 11 1736 45
rect 1770 11 1781 45
rect 1725 -23 1781 11
rect 1725 -57 1736 -23
rect 1770 -57 1781 -23
rect 1725 -91 1781 -57
rect 1725 -125 1736 -91
rect 1770 -125 1781 -91
rect 1725 -159 1781 -125
rect 1725 -193 1736 -159
rect 1770 -193 1781 -159
rect 1725 -205 1781 -193
rect 1941 725 1997 795
rect 1941 691 1952 725
rect 1986 691 1997 725
rect 1941 657 1997 691
rect 1941 623 1952 657
rect 1986 623 1997 657
rect 1941 589 1997 623
rect 1941 555 1952 589
rect 1986 555 1997 589
rect 1941 521 1997 555
rect 1941 487 1952 521
rect 1986 487 1997 521
rect 1941 453 1997 487
rect 1941 419 1952 453
rect 1986 419 1997 453
rect 1941 385 1997 419
rect 1941 351 1952 385
rect 1986 351 1997 385
rect 1941 317 1997 351
rect 1941 283 1952 317
rect 1986 283 1997 317
rect 1941 249 1997 283
rect 1941 215 1952 249
rect 1986 215 1997 249
rect 1941 181 1997 215
rect 1941 147 1952 181
rect 1986 147 1997 181
rect 1941 113 1997 147
rect 1941 79 1952 113
rect 1986 79 1997 113
rect 1941 45 1997 79
rect 1941 11 1952 45
rect 1986 11 1997 45
rect 1941 -23 1997 11
rect 1941 -57 1952 -23
rect 1986 -57 1997 -23
rect 1941 -91 1997 -57
rect 1941 -125 1952 -91
rect 1986 -125 1997 -91
rect 1941 -159 1997 -125
rect 1941 -193 1952 -159
rect 1986 -193 1997 -159
rect 1941 -205 1997 -193
rect 2157 725 2210 795
rect 2157 691 2168 725
rect 2202 691 2210 725
rect 2157 657 2210 691
rect 2157 623 2168 657
rect 2202 623 2210 657
rect 2157 589 2210 623
rect 2157 555 2168 589
rect 2202 555 2210 589
rect 2157 521 2210 555
rect 2157 487 2168 521
rect 2202 487 2210 521
rect 2157 453 2210 487
rect 2157 419 2168 453
rect 2202 419 2210 453
rect 2157 385 2210 419
rect 2157 351 2168 385
rect 2202 351 2210 385
rect 2157 317 2210 351
rect 2157 283 2168 317
rect 2202 283 2210 317
rect 2157 249 2210 283
rect 2157 215 2168 249
rect 2202 215 2210 249
rect 2157 181 2210 215
rect 2157 147 2168 181
rect 2202 147 2210 181
rect 2157 113 2210 147
rect 2157 79 2168 113
rect 2202 79 2210 113
rect 2157 45 2210 79
rect 2157 11 2168 45
rect 2202 11 2210 45
rect 2157 -23 2210 11
rect 2157 -57 2168 -23
rect 2202 -57 2210 -23
rect 2157 -91 2210 -57
rect 2157 -125 2168 -91
rect 2202 -125 2210 -91
rect 2157 -159 2210 -125
rect 2157 -193 2168 -159
rect 2202 -193 2210 -159
rect 2157 -205 2210 -193
rect 2270 725 2323 795
rect 2270 691 2278 725
rect 2312 691 2323 725
rect 2270 657 2323 691
rect 2270 623 2278 657
rect 2312 623 2323 657
rect 2270 589 2323 623
rect 2270 555 2278 589
rect 2312 555 2323 589
rect 2270 521 2323 555
rect 2270 487 2278 521
rect 2312 487 2323 521
rect 2270 453 2323 487
rect 2270 419 2278 453
rect 2312 419 2323 453
rect 2270 385 2323 419
rect 2270 351 2278 385
rect 2312 351 2323 385
rect 2270 317 2323 351
rect 2270 283 2278 317
rect 2312 283 2323 317
rect 2270 249 2323 283
rect 2270 215 2278 249
rect 2312 215 2323 249
rect 2270 181 2323 215
rect 2270 147 2278 181
rect 2312 147 2323 181
rect 2270 113 2323 147
rect 2270 79 2278 113
rect 2312 79 2323 113
rect 2270 45 2323 79
rect 2270 11 2278 45
rect 2312 11 2323 45
rect 2270 -23 2323 11
rect 2270 -57 2278 -23
rect 2312 -57 2323 -23
rect 2270 -91 2323 -57
rect 2270 -125 2278 -91
rect 2312 -125 2323 -91
rect 2270 -159 2323 -125
rect 2270 -193 2278 -159
rect 2312 -193 2323 -159
rect 2270 -205 2323 -193
rect 2483 725 2536 795
rect 2483 691 2494 725
rect 2528 691 2536 725
rect 2483 657 2536 691
rect 2483 623 2494 657
rect 2528 623 2536 657
rect 2483 589 2536 623
rect 2483 555 2494 589
rect 2528 555 2536 589
rect 2483 521 2536 555
rect 2483 487 2494 521
rect 2528 487 2536 521
rect 2483 453 2536 487
rect 2483 419 2494 453
rect 2528 419 2536 453
rect 2483 385 2536 419
rect 2483 351 2494 385
rect 2528 351 2536 385
rect 2483 317 2536 351
rect 2483 283 2494 317
rect 2528 283 2536 317
rect 2483 249 2536 283
rect 2483 215 2494 249
rect 2528 215 2536 249
rect 2483 181 2536 215
rect 2483 147 2494 181
rect 2528 147 2536 181
rect 2483 113 2536 147
rect 2483 79 2494 113
rect 2528 79 2536 113
rect 2483 45 2536 79
rect 2483 11 2494 45
rect 2528 11 2536 45
rect 2483 -23 2536 11
rect 2483 -57 2494 -23
rect 2528 -57 2536 -23
rect 2483 -91 2536 -57
rect 2483 -125 2494 -91
rect 2528 -125 2536 -91
rect 2483 -159 2536 -125
rect 2483 -193 2494 -159
rect 2528 -193 2536 -159
rect 2483 -205 2536 -193
<< mvpdiff >>
rect 642 2002 1642 2010
rect 642 1968 654 2002
rect 688 1968 722 2002
rect 756 1968 790 2002
rect 824 1968 858 2002
rect 892 1968 926 2002
rect 960 1968 994 2002
rect 1028 1968 1062 2002
rect 1096 1968 1130 2002
rect 1164 1968 1198 2002
rect 1232 1968 1266 2002
rect 1300 1968 1334 2002
rect 1368 1968 1402 2002
rect 1436 1968 1470 2002
rect 1504 1968 1538 2002
rect 1572 1968 1642 2002
rect 642 1957 1642 1968
rect 642 1786 1642 1797
rect 642 1752 654 1786
rect 688 1752 722 1786
rect 756 1752 790 1786
rect 824 1752 858 1786
rect 892 1752 926 1786
rect 960 1752 994 1786
rect 1028 1752 1062 1786
rect 1096 1752 1130 1786
rect 1164 1752 1198 1786
rect 1232 1752 1266 1786
rect 1300 1752 1334 1786
rect 1368 1752 1402 1786
rect 1436 1752 1470 1786
rect 1504 1752 1538 1786
rect 1572 1752 1642 1786
rect 642 1741 1642 1752
rect 642 1570 1642 1581
rect 642 1536 654 1570
rect 688 1536 722 1570
rect 756 1536 790 1570
rect 824 1536 858 1570
rect 892 1536 926 1570
rect 960 1536 994 1570
rect 1028 1536 1062 1570
rect 1096 1536 1130 1570
rect 1164 1536 1198 1570
rect 1232 1536 1266 1570
rect 1300 1536 1334 1570
rect 1368 1536 1402 1570
rect 1436 1536 1470 1570
rect 1504 1536 1538 1570
rect 1572 1536 1642 1570
rect 642 1528 1642 1536
<< ndiffc >>
rect 210 27 244 61
rect 210 -41 244 -7
rect 210 -109 244 -75
rect 316 27 350 61
rect 316 -41 350 -7
rect 316 -109 350 -75
rect 422 27 456 61
rect 422 -41 456 -7
rect 422 -109 456 -75
rect 528 27 562 61
rect 528 -41 562 -7
rect 528 -109 562 -75
rect 638 27 672 61
rect 638 -41 672 -7
rect 638 -109 672 -75
rect 744 27 778 61
rect 744 -41 778 -7
rect 744 -109 778 -75
rect 850 27 884 61
rect 850 -41 884 -7
rect 850 -109 884 -75
rect 956 27 990 61
rect 956 -41 990 -7
rect 956 -109 990 -75
rect 1062 27 1096 61
rect 1062 -41 1096 -7
rect 1062 -109 1096 -75
rect 1168 27 1202 61
rect 1168 -41 1202 -7
rect 1168 -109 1202 -75
<< pdiffc >>
rect 1430 3552 1464 3586
rect 1498 3552 1532 3586
rect 1566 3552 1600 3586
rect 690 3446 724 3480
rect 758 3446 792 3480
rect 826 3446 860 3480
rect 894 3446 928 3480
rect 962 3446 996 3480
rect 1030 3446 1064 3480
rect 1098 3446 1132 3480
rect 1166 3446 1200 3480
rect 1430 3446 1464 3480
rect 1498 3446 1532 3480
rect 1566 3446 1600 3480
rect 690 3340 724 3374
rect 758 3340 792 3374
rect 826 3340 860 3374
rect 894 3340 928 3374
rect 962 3340 996 3374
rect 1030 3340 1064 3374
rect 1098 3340 1132 3374
rect 1166 3340 1200 3374
rect 1430 3340 1464 3374
rect 1498 3340 1532 3374
rect 1566 3340 1600 3374
rect 682 3230 716 3264
rect 750 3230 784 3264
rect 818 3230 852 3264
rect 886 3230 920 3264
rect 954 3230 988 3264
rect 1022 3230 1056 3264
rect 1090 3230 1124 3264
rect 1158 3230 1192 3264
rect 1226 3230 1260 3264
rect 1294 3230 1328 3264
rect 1362 3230 1396 3264
rect 1430 3230 1464 3264
rect 1498 3230 1532 3264
rect 1566 3230 1600 3264
rect 682 3124 716 3158
rect 750 3124 784 3158
rect 818 3124 852 3158
rect 886 3124 920 3158
rect 954 3124 988 3158
rect 1022 3124 1056 3158
rect 1090 3124 1124 3158
rect 1158 3124 1192 3158
rect 1226 3124 1260 3158
rect 1294 3124 1328 3158
rect 1362 3124 1396 3158
rect 1430 3124 1464 3158
rect 1498 3124 1532 3158
rect 1566 3124 1600 3158
rect 682 3018 716 3052
rect 750 3018 784 3052
rect 818 3018 852 3052
rect 886 3018 920 3052
rect 954 3018 988 3052
rect 1022 3018 1056 3052
rect 1090 3018 1124 3052
rect 1158 3018 1192 3052
rect 1226 3018 1260 3052
rect 1294 3018 1328 3052
rect 1362 3018 1396 3052
rect 1430 3018 1464 3052
rect 1498 3018 1532 3052
rect 1566 3018 1600 3052
rect 682 2908 716 2942
rect 750 2908 784 2942
rect 818 2908 852 2942
rect 886 2908 920 2942
rect 954 2908 988 2942
rect 1022 2908 1056 2942
rect 1090 2908 1124 2942
rect 1158 2908 1192 2942
rect 1226 2908 1260 2942
rect 1294 2908 1328 2942
rect 1362 2908 1396 2942
rect 1430 2908 1464 2942
rect 1498 2908 1532 2942
rect 1566 2908 1600 2942
rect 682 2802 716 2836
rect 750 2802 784 2836
rect 818 2802 852 2836
rect 886 2802 920 2836
rect 954 2802 988 2836
rect 1022 2802 1056 2836
rect 1090 2802 1124 2836
rect 1158 2802 1192 2836
rect 1226 2802 1260 2836
rect 1294 2802 1328 2836
rect 1362 2802 1396 2836
rect 1430 2802 1464 2836
rect 1498 2802 1532 2836
rect 1566 2802 1600 2836
rect 682 2696 716 2730
rect 750 2696 784 2730
rect 818 2696 852 2730
rect 886 2696 920 2730
rect 954 2696 988 2730
rect 1022 2696 1056 2730
rect 1090 2696 1124 2730
rect 1158 2696 1192 2730
rect 1226 2696 1260 2730
rect 1294 2696 1328 2730
rect 1362 2696 1396 2730
rect 1430 2696 1464 2730
rect 1498 2696 1532 2730
rect 1566 2696 1600 2730
rect 682 2590 716 2624
rect 750 2590 784 2624
rect 818 2590 852 2624
rect 886 2590 920 2624
rect 954 2590 988 2624
rect 1022 2590 1056 2624
rect 1090 2590 1124 2624
rect 1158 2590 1192 2624
rect 1226 2590 1260 2624
rect 1294 2590 1328 2624
rect 1362 2590 1396 2624
rect 1430 2590 1464 2624
rect 1498 2590 1532 2624
rect 1566 2590 1600 2624
rect 682 2484 716 2518
rect 750 2484 784 2518
rect 818 2484 852 2518
rect 886 2484 920 2518
rect 954 2484 988 2518
rect 1022 2484 1056 2518
rect 1090 2484 1124 2518
rect 1158 2484 1192 2518
rect 1226 2484 1260 2518
rect 1294 2484 1328 2518
rect 1362 2484 1396 2518
rect 1430 2484 1464 2518
rect 1498 2484 1532 2518
rect 1566 2484 1600 2518
<< mvndiffc >>
rect 220 743 254 777
rect 220 675 254 709
rect 220 607 254 641
rect 436 743 470 777
rect 436 675 470 709
rect 436 607 470 641
rect 546 743 580 777
rect 546 675 580 709
rect 546 607 580 641
rect 762 743 796 777
rect 762 675 796 709
rect 762 607 796 641
rect 978 743 1012 777
rect 978 675 1012 709
rect 978 607 1012 641
rect 1194 743 1228 777
rect 1194 675 1228 709
rect 1194 607 1228 641
rect 1304 691 1338 725
rect 1304 623 1338 657
rect 1304 555 1338 589
rect 1304 487 1338 521
rect 1304 419 1338 453
rect 1304 351 1338 385
rect 1304 283 1338 317
rect 1304 215 1338 249
rect 1304 147 1338 181
rect 1304 79 1338 113
rect 1304 11 1338 45
rect 1304 -57 1338 -23
rect 1304 -125 1338 -91
rect 1304 -193 1338 -159
rect 1520 691 1554 725
rect 1520 623 1554 657
rect 1520 555 1554 589
rect 1520 487 1554 521
rect 1520 419 1554 453
rect 1520 351 1554 385
rect 1520 283 1554 317
rect 1520 215 1554 249
rect 1520 147 1554 181
rect 1520 79 1554 113
rect 1520 11 1554 45
rect 1520 -57 1554 -23
rect 1520 -125 1554 -91
rect 1520 -193 1554 -159
rect 1736 691 1770 725
rect 1736 623 1770 657
rect 1736 555 1770 589
rect 1736 487 1770 521
rect 1736 419 1770 453
rect 1736 351 1770 385
rect 1736 283 1770 317
rect 1736 215 1770 249
rect 1736 147 1770 181
rect 1736 79 1770 113
rect 1736 11 1770 45
rect 1736 -57 1770 -23
rect 1736 -125 1770 -91
rect 1736 -193 1770 -159
rect 1952 691 1986 725
rect 1952 623 1986 657
rect 1952 555 1986 589
rect 1952 487 1986 521
rect 1952 419 1986 453
rect 1952 351 1986 385
rect 1952 283 1986 317
rect 1952 215 1986 249
rect 1952 147 1986 181
rect 1952 79 1986 113
rect 1952 11 1986 45
rect 1952 -57 1986 -23
rect 1952 -125 1986 -91
rect 1952 -193 1986 -159
rect 2168 691 2202 725
rect 2168 623 2202 657
rect 2168 555 2202 589
rect 2168 487 2202 521
rect 2168 419 2202 453
rect 2168 351 2202 385
rect 2168 283 2202 317
rect 2168 215 2202 249
rect 2168 147 2202 181
rect 2168 79 2202 113
rect 2168 11 2202 45
rect 2168 -57 2202 -23
rect 2168 -125 2202 -91
rect 2168 -193 2202 -159
rect 2278 691 2312 725
rect 2278 623 2312 657
rect 2278 555 2312 589
rect 2278 487 2312 521
rect 2278 419 2312 453
rect 2278 351 2312 385
rect 2278 283 2312 317
rect 2278 215 2312 249
rect 2278 147 2312 181
rect 2278 79 2312 113
rect 2278 11 2312 45
rect 2278 -57 2312 -23
rect 2278 -125 2312 -91
rect 2278 -193 2312 -159
rect 2494 691 2528 725
rect 2494 623 2528 657
rect 2494 555 2528 589
rect 2494 487 2528 521
rect 2494 419 2528 453
rect 2494 351 2528 385
rect 2494 283 2528 317
rect 2494 215 2528 249
rect 2494 147 2528 181
rect 2494 79 2528 113
rect 2494 11 2528 45
rect 2494 -57 2528 -23
rect 2494 -125 2528 -91
rect 2494 -193 2528 -159
<< mvpdiffc >>
rect 654 1968 688 2002
rect 722 1968 756 2002
rect 790 1968 824 2002
rect 858 1968 892 2002
rect 926 1968 960 2002
rect 994 1968 1028 2002
rect 1062 1968 1096 2002
rect 1130 1968 1164 2002
rect 1198 1968 1232 2002
rect 1266 1968 1300 2002
rect 1334 1968 1368 2002
rect 1402 1968 1436 2002
rect 1470 1968 1504 2002
rect 1538 1968 1572 2002
rect 654 1752 688 1786
rect 722 1752 756 1786
rect 790 1752 824 1786
rect 858 1752 892 1786
rect 926 1752 960 1786
rect 994 1752 1028 1786
rect 1062 1752 1096 1786
rect 1130 1752 1164 1786
rect 1198 1752 1232 1786
rect 1266 1752 1300 1786
rect 1334 1752 1368 1786
rect 1402 1752 1436 1786
rect 1470 1752 1504 1786
rect 1538 1752 1572 1786
rect 654 1536 688 1570
rect 722 1536 756 1570
rect 790 1536 824 1570
rect 858 1536 892 1570
rect 926 1536 960 1570
rect 994 1536 1028 1570
rect 1062 1536 1096 1570
rect 1130 1536 1164 1570
rect 1198 1536 1232 1570
rect 1266 1536 1300 1570
rect 1334 1536 1368 1570
rect 1402 1536 1436 1570
rect 1470 1536 1504 1570
rect 1538 1536 1572 1570
<< nsubdiff >>
rect 643 3544 677 3578
rect 711 3544 745 3578
rect 779 3544 813 3578
rect 847 3544 881 3578
rect 915 3544 949 3578
rect 983 3544 1017 3578
rect 1051 3544 1085 3578
rect 1119 3544 1181 3578
rect 1694 3514 1728 3563
rect 1694 3446 1728 3480
rect 1694 3378 1728 3412
rect 1694 3310 1728 3344
rect 1694 3242 1728 3276
rect 1694 3174 1728 3208
rect 1694 3106 1728 3140
rect 1694 3038 1728 3072
rect 1694 2970 1728 3004
rect 1694 2902 1728 2936
rect 1694 2834 1728 2868
rect 1694 2766 1728 2800
rect 1694 2698 1728 2732
rect 1694 2630 1728 2664
<< mvpsubdiff >>
rect 230 441 254 475
rect 288 441 324 475
rect 358 441 393 475
rect 427 441 462 475
rect 496 441 531 475
rect 565 441 600 475
rect 634 441 669 475
rect 703 441 738 475
rect 772 441 807 475
rect 841 441 876 475
rect 910 441 945 475
rect 979 441 1014 475
rect 1048 441 1083 475
rect 1117 441 1152 475
rect 1186 441 1210 475
rect 172 -315 196 -281
rect 230 -315 267 -281
rect 301 -315 338 -281
rect 372 -315 408 -281
rect 442 -315 478 -281
rect 512 -315 548 -281
rect 582 -315 618 -281
rect 652 -315 688 -281
rect 722 -315 758 -281
rect 792 -315 828 -281
rect 862 -315 898 -281
rect 932 -315 968 -281
rect 1002 -315 1038 -281
rect 1072 -315 1108 -281
rect 1142 -315 1178 -281
rect 1212 -315 1248 -281
rect 1282 -315 1318 -281
rect 1352 -315 1388 -281
rect 1422 -315 1458 -281
rect 1492 -315 1528 -281
rect 1562 -315 1598 -281
rect 1632 -315 1668 -281
rect 1702 -315 1738 -281
rect 1772 -315 1808 -281
rect 1842 -315 1878 -281
rect 1912 -315 1948 -281
rect 1982 -315 2018 -281
rect 2052 -315 2088 -281
rect 2122 -315 2158 -281
rect 2192 -315 2228 -281
rect 2262 -315 2298 -281
rect 2332 -315 2368 -281
rect 2402 -315 2438 -281
rect 2472 -315 2496 -281
<< mvnsubdiff >>
rect 1716 1937 1750 2009
rect 1716 1869 1750 1903
rect 1716 1801 1750 1835
rect 1716 1733 1750 1767
rect 1716 1665 1750 1699
rect 1716 1597 1750 1631
rect 1716 1529 1750 1563
<< nsubdiffcont >>
rect 677 3544 711 3578
rect 745 3544 779 3578
rect 813 3544 847 3578
rect 881 3544 915 3578
rect 949 3544 983 3578
rect 1017 3544 1051 3578
rect 1085 3544 1119 3578
rect 1694 3480 1728 3514
rect 1694 3412 1728 3446
rect 1694 3344 1728 3378
rect 1694 3276 1728 3310
rect 1694 3208 1728 3242
rect 1694 3140 1728 3174
rect 1694 3072 1728 3106
rect 1694 3004 1728 3038
rect 1694 2936 1728 2970
rect 1694 2868 1728 2902
rect 1694 2800 1728 2834
rect 1694 2732 1728 2766
rect 1694 2664 1728 2698
<< mvpsubdiffcont >>
rect 254 441 288 475
rect 324 441 358 475
rect 393 441 427 475
rect 462 441 496 475
rect 531 441 565 475
rect 600 441 634 475
rect 669 441 703 475
rect 738 441 772 475
rect 807 441 841 475
rect 876 441 910 475
rect 945 441 979 475
rect 1014 441 1048 475
rect 1083 441 1117 475
rect 1152 441 1186 475
rect 196 -315 230 -281
rect 267 -315 301 -281
rect 338 -315 372 -281
rect 408 -315 442 -281
rect 478 -315 512 -281
rect 548 -315 582 -281
rect 618 -315 652 -281
rect 688 -315 722 -281
rect 758 -315 792 -281
rect 828 -315 862 -281
rect 898 -315 932 -281
rect 968 -315 1002 -281
rect 1038 -315 1072 -281
rect 1108 -315 1142 -281
rect 1178 -315 1212 -281
rect 1248 -315 1282 -281
rect 1318 -315 1352 -281
rect 1388 -315 1422 -281
rect 1458 -315 1492 -281
rect 1528 -315 1562 -281
rect 1598 -315 1632 -281
rect 1668 -315 1702 -281
rect 1738 -315 1772 -281
rect 1808 -315 1842 -281
rect 1878 -315 1912 -281
rect 1948 -315 1982 -281
rect 2018 -315 2052 -281
rect 2088 -315 2122 -281
rect 2158 -315 2192 -281
rect 2228 -315 2262 -281
rect 2298 -315 2332 -281
rect 2368 -315 2402 -281
rect 2438 -315 2472 -281
<< mvnsubdiffcont >>
rect 1716 1903 1750 1937
rect 1716 1835 1750 1869
rect 1716 1767 1750 1801
rect 1716 1699 1750 1733
rect 1716 1631 1750 1665
rect 1716 1563 1750 1597
<< poly >>
rect 1314 3525 1412 3541
rect 1314 3491 1330 3525
rect 1364 3491 1412 3525
rect 1612 3491 1644 3541
rect 446 3435 580 3441
rect 1314 3435 1380 3491
rect 446 3425 612 3435
rect 446 3391 462 3425
rect 496 3391 530 3425
rect 564 3391 612 3425
rect 446 3385 612 3391
rect 1212 3385 1244 3435
rect 1314 3401 1330 3435
rect 1364 3401 1412 3435
rect 1314 3385 1412 3401
rect 1612 3385 1644 3435
rect 446 3375 580 3385
rect 446 3219 580 3235
rect 446 3185 462 3219
rect 496 3185 530 3219
rect 564 3185 612 3219
rect 446 3169 612 3185
rect 1612 3169 1644 3219
rect 446 3113 580 3121
rect 446 3105 612 3113
rect 446 3071 462 3105
rect 496 3071 530 3105
rect 564 3071 612 3105
rect 446 3063 612 3071
rect 1612 3063 1644 3113
rect 446 3055 580 3063
rect 446 2897 580 2907
rect 446 2891 612 2897
rect 446 2857 462 2891
rect 496 2857 530 2891
rect 564 2857 612 2891
rect 446 2847 612 2857
rect 1612 2847 1644 2897
rect 446 2841 580 2847
rect 514 2775 612 2791
rect 514 2741 530 2775
rect 564 2741 612 2775
rect 1612 2741 1644 2791
rect 514 2685 580 2741
rect 514 2677 612 2685
rect 514 2643 530 2677
rect 564 2643 612 2677
rect 514 2635 612 2643
rect 1612 2635 1644 2685
rect 514 2579 580 2635
rect 514 2545 530 2579
rect 564 2545 612 2579
rect 514 2529 612 2545
rect 1612 2529 1644 2579
rect 544 1941 642 1957
rect 544 1907 560 1941
rect 594 1907 642 1941
rect 544 1864 642 1907
rect 544 1830 560 1864
rect 594 1830 642 1864
rect 544 1797 642 1830
rect 1642 1797 1674 1957
rect 544 1787 610 1797
rect 544 1753 560 1787
rect 594 1753 610 1787
rect 544 1741 610 1753
rect 544 1709 642 1741
rect 544 1675 560 1709
rect 594 1675 642 1709
rect 544 1631 642 1675
rect 544 1597 560 1631
rect 594 1597 642 1631
rect 544 1581 642 1597
rect 1642 1581 1674 1741
rect 265 877 425 893
rect 265 843 281 877
rect 315 843 375 877
rect 409 843 425 877
rect 265 795 425 843
rect 591 877 1183 893
rect 591 843 607 877
rect 641 843 683 877
rect 717 843 758 877
rect 792 843 833 877
rect 867 843 908 877
rect 942 843 983 877
rect 1017 843 1058 877
rect 1092 843 1133 877
rect 1167 843 1183 877
rect 591 827 1183 843
rect 591 795 751 827
rect 807 795 967 827
rect 1023 795 1183 827
rect 1349 877 2157 893
rect 1349 843 1365 877
rect 1399 843 1440 877
rect 1474 843 1515 877
rect 1549 843 1589 877
rect 1623 843 1663 877
rect 1697 843 1737 877
rect 1771 843 1811 877
rect 1845 843 1885 877
rect 1919 843 1959 877
rect 1993 843 2033 877
rect 2067 843 2107 877
rect 2141 843 2157 877
rect 1349 827 2157 843
rect 1349 795 1509 827
rect 1565 795 1725 827
rect 1781 795 1941 827
rect 1997 795 2157 827
rect 2323 877 2483 893
rect 2323 843 2339 877
rect 2373 843 2433 877
rect 2467 843 2483 877
rect 2323 795 2483 843
rect 265 563 425 595
rect 591 563 751 595
rect 807 563 967 595
rect 1023 563 1183 595
rect 255 155 517 171
rect 255 121 271 155
rect 305 121 369 155
rect 403 121 467 155
rect 501 121 517 155
rect 255 105 517 121
rect 577 155 733 171
rect 577 121 593 155
rect 627 121 683 155
rect 717 121 733 155
rect 577 105 733 121
rect 255 73 305 105
rect 361 73 411 105
rect 467 73 517 105
rect 683 73 733 105
rect 789 155 945 171
rect 789 121 805 155
rect 839 121 895 155
rect 929 121 945 155
rect 789 105 945 121
rect 789 73 839 105
rect 895 73 945 105
rect 1001 155 1157 171
rect 1001 121 1017 155
rect 1051 121 1107 155
rect 1141 121 1157 155
rect 1001 105 1157 121
rect 1001 73 1051 105
rect 1107 73 1157 105
rect 255 -159 305 -127
rect 361 -159 411 -127
rect 467 -159 517 -127
rect 683 -159 733 -127
rect 789 -159 839 -127
rect 895 -159 945 -127
rect 1001 -159 1051 -127
rect 1107 -159 1157 -127
rect 1349 -237 1509 -205
rect 1565 -237 1725 -205
rect 1781 -237 1941 -205
rect 1997 -237 2157 -205
rect 2323 -237 2483 -205
<< polycont >>
rect 1330 3491 1364 3525
rect 462 3391 496 3425
rect 530 3391 564 3425
rect 1330 3401 1364 3435
rect 462 3185 496 3219
rect 530 3185 564 3219
rect 462 3071 496 3105
rect 530 3071 564 3105
rect 462 2857 496 2891
rect 530 2857 564 2891
rect 530 2741 564 2775
rect 530 2643 564 2677
rect 530 2545 564 2579
rect 560 1907 594 1941
rect 560 1830 594 1864
rect 560 1753 594 1787
rect 560 1675 594 1709
rect 560 1597 594 1631
rect 281 843 315 877
rect 375 843 409 877
rect 607 843 641 877
rect 683 843 717 877
rect 758 843 792 877
rect 833 843 867 877
rect 908 843 942 877
rect 983 843 1017 877
rect 1058 843 1092 877
rect 1133 843 1167 877
rect 1365 843 1399 877
rect 1440 843 1474 877
rect 1515 843 1549 877
rect 1589 843 1623 877
rect 1663 843 1697 877
rect 1737 843 1771 877
rect 1811 843 1845 877
rect 1885 843 1919 877
rect 1959 843 1993 877
rect 2033 843 2067 877
rect 2107 843 2141 877
rect 2339 843 2373 877
rect 2433 843 2467 877
rect 271 121 305 155
rect 369 121 403 155
rect 467 121 501 155
rect 593 121 627 155
rect 683 121 717 155
rect 805 121 839 155
rect 895 121 929 155
rect 1017 121 1051 155
rect 1107 121 1141 155
<< locali >>
rect 643 3544 673 3578
rect 711 3544 745 3578
rect 784 3544 813 3578
rect 861 3544 881 3578
rect 938 3544 949 3578
rect 1015 3544 1017 3578
rect 1051 3544 1058 3578
rect 1119 3544 1135 3578
rect 1169 3544 1181 3578
rect 1414 3552 1430 3586
rect 1464 3552 1494 3586
rect 1532 3552 1566 3586
rect 1600 3552 1616 3586
rect 1330 3526 1364 3541
rect 724 3446 757 3480
rect 792 3446 826 3480
rect 874 3446 894 3480
rect 956 3446 962 3480
rect 996 3446 1004 3480
rect 1064 3446 1086 3480
rect 1132 3446 1166 3480
rect 1202 3446 1216 3480
rect 1330 3454 1364 3491
rect 1694 3534 1728 3563
rect 1464 3446 1486 3480
rect 1532 3446 1566 3480
rect 1600 3446 1616 3480
rect 1694 3462 1728 3480
rect 446 3391 452 3425
rect 496 3391 524 3425
rect 564 3391 580 3425
rect 1330 3385 1364 3401
rect 1694 3390 1728 3412
rect 674 3340 690 3374
rect 724 3340 746 3374
rect 792 3340 826 3374
rect 865 3340 894 3374
rect 950 3340 962 3374
rect 996 3340 1001 3374
rect 1064 3340 1086 3374
rect 1132 3340 1166 3374
rect 1204 3340 1216 3374
rect 1414 3340 1430 3374
rect 1464 3340 1494 3374
rect 1532 3340 1566 3374
rect 1600 3340 1616 3374
rect 1694 3318 1728 3344
rect 716 3230 745 3264
rect 784 3230 818 3264
rect 858 3230 886 3264
rect 937 3230 954 3264
rect 1016 3230 1022 3264
rect 1056 3230 1061 3264
rect 1124 3230 1140 3264
rect 1192 3230 1219 3264
rect 1260 3230 1294 3264
rect 1331 3230 1362 3264
rect 1409 3230 1430 3264
rect 1487 3230 1498 3264
rect 1532 3230 1566 3264
rect 1600 3230 1616 3264
rect 1694 3246 1728 3276
rect 446 3212 462 3219
rect 496 3212 530 3219
rect 446 3185 454 3212
rect 496 3185 526 3212
rect 564 3185 580 3219
rect 488 3178 526 3185
rect 1694 3174 1728 3208
rect 666 3124 682 3158
rect 716 3124 750 3158
rect 784 3124 795 3158
rect 852 3124 874 3158
rect 920 3124 953 3158
rect 988 3124 1022 3158
rect 1066 3124 1090 3158
rect 1145 3124 1158 3158
rect 1224 3124 1226 3158
rect 1260 3124 1269 3158
rect 1328 3124 1348 3158
rect 1396 3124 1426 3158
rect 1464 3124 1498 3158
rect 1538 3124 1566 3158
rect 1694 3106 1728 3140
rect 446 3071 450 3105
rect 496 3071 522 3105
rect 564 3071 580 3105
rect 716 3018 745 3052
rect 784 3018 818 3052
rect 858 3018 886 3052
rect 937 3018 954 3052
rect 1016 3018 1022 3052
rect 1056 3018 1061 3052
rect 1124 3018 1140 3052
rect 1192 3018 1219 3052
rect 1260 3018 1294 3052
rect 1331 3018 1362 3052
rect 1409 3018 1430 3052
rect 1487 3018 1498 3052
rect 1532 3018 1566 3052
rect 1600 3018 1616 3052
rect 1694 3038 1728 3068
rect 1694 2970 1728 2995
rect 716 2908 745 2942
rect 784 2908 818 2942
rect 858 2908 886 2942
rect 937 2908 954 2942
rect 1016 2908 1022 2942
rect 1056 2908 1061 2942
rect 1124 2908 1140 2942
rect 1192 2908 1219 2942
rect 1260 2908 1294 2942
rect 1331 2908 1362 2942
rect 1409 2908 1430 2942
rect 1487 2908 1498 2942
rect 1532 2908 1566 2942
rect 1600 2908 1616 2942
rect 1694 2902 1728 2922
rect 446 2857 452 2891
rect 496 2857 524 2891
rect 564 2857 580 2891
rect 666 2802 682 2836
rect 716 2802 750 2836
rect 784 2802 795 2836
rect 852 2802 874 2836
rect 920 2802 953 2836
rect 988 2802 1022 2836
rect 1066 2802 1090 2836
rect 1145 2802 1158 2836
rect 1224 2802 1226 2836
rect 1260 2802 1269 2836
rect 1328 2802 1348 2836
rect 1396 2802 1426 2836
rect 1464 2802 1498 2836
rect 1538 2802 1566 2836
rect 1694 2834 1728 2849
rect 530 2775 564 2791
rect 530 2683 564 2731
rect 1694 2766 1728 2776
rect 716 2696 745 2730
rect 784 2696 818 2730
rect 858 2696 886 2730
rect 937 2696 954 2730
rect 1016 2696 1022 2730
rect 1056 2696 1061 2730
rect 1124 2696 1140 2730
rect 1192 2696 1219 2730
rect 1260 2696 1294 2730
rect 1331 2696 1362 2730
rect 1409 2696 1430 2730
rect 1487 2696 1498 2730
rect 1532 2696 1566 2730
rect 1600 2696 1616 2730
rect 1694 2698 1728 2703
rect 530 2601 564 2643
rect 666 2590 682 2624
rect 716 2590 750 2624
rect 784 2590 795 2624
rect 852 2590 874 2624
rect 920 2590 953 2624
rect 988 2590 1022 2624
rect 1066 2590 1090 2624
rect 1145 2590 1158 2624
rect 1224 2590 1226 2624
rect 1260 2590 1269 2624
rect 1328 2590 1348 2624
rect 1396 2590 1426 2624
rect 1464 2590 1498 2624
rect 1538 2590 1566 2624
rect 530 2529 564 2545
rect 716 2484 745 2518
rect 784 2484 818 2518
rect 858 2484 886 2518
rect 937 2484 954 2518
rect 1016 2484 1022 2518
rect 1056 2484 1061 2518
rect 1124 2484 1140 2518
rect 1192 2484 1219 2518
rect 1260 2484 1294 2518
rect 1331 2484 1362 2518
rect 1409 2484 1430 2518
rect 1487 2484 1498 2518
rect 1532 2484 1566 2518
rect 1600 2484 1616 2518
rect 638 1968 654 2002
rect 688 1968 699 2002
rect 756 1968 776 2002
rect 824 1968 853 2002
rect 892 1968 926 2002
rect 964 1968 994 2002
rect 1041 1968 1062 2002
rect 1118 1968 1130 2002
rect 1195 1968 1198 2002
rect 1232 1968 1238 2002
rect 1300 1968 1314 2002
rect 1368 1968 1390 2002
rect 1436 1968 1466 2002
rect 1504 1968 1538 2002
rect 1576 1968 1588 2002
rect 1716 1997 1750 2009
rect 560 1941 594 1957
rect 560 1864 594 1881
rect 560 1823 594 1830
rect 560 1787 594 1789
rect 1716 1937 1750 1963
rect 1716 1869 1750 1891
rect 1716 1801 1750 1819
rect 560 1731 594 1753
rect 638 1752 654 1786
rect 688 1752 699 1786
rect 756 1752 777 1786
rect 824 1752 855 1786
rect 892 1752 926 1786
rect 967 1752 994 1786
rect 1045 1752 1062 1786
rect 1123 1752 1130 1786
rect 1164 1752 1167 1786
rect 1232 1752 1245 1786
rect 1300 1752 1322 1786
rect 1368 1752 1399 1786
rect 1436 1752 1470 1786
rect 1510 1752 1538 1786
rect 1587 1752 1588 1786
rect 560 1638 594 1675
rect 560 1581 594 1597
rect 1716 1733 1750 1747
rect 1716 1665 1750 1675
rect 1716 1597 1750 1602
rect 638 1536 654 1570
rect 688 1536 699 1570
rect 756 1536 777 1570
rect 824 1536 855 1570
rect 892 1536 926 1570
rect 967 1536 994 1570
rect 1045 1536 1062 1570
rect 1123 1536 1130 1570
rect 1164 1536 1167 1570
rect 1232 1536 1245 1570
rect 1300 1536 1322 1570
rect 1368 1536 1399 1570
rect 1436 1536 1470 1570
rect 1510 1536 1538 1570
rect 1587 1536 1588 1570
rect 265 843 281 877
rect 325 843 363 877
rect 409 843 425 877
rect 591 843 607 877
rect 665 843 683 877
rect 745 843 758 877
rect 825 843 833 877
rect 867 843 871 877
rect 905 843 908 877
rect 942 843 950 877
rect 1017 843 1029 877
rect 1092 843 1108 877
rect 1167 843 1183 877
rect 1349 843 1365 877
rect 1403 843 1440 877
rect 1478 843 1515 877
rect 1553 843 1589 877
rect 1628 843 1663 877
rect 1702 843 1737 877
rect 1776 843 1811 877
rect 1850 843 1885 877
rect 1924 843 1959 877
rect 1998 843 2033 877
rect 2072 843 2107 877
rect 2146 843 2157 877
rect 2323 843 2339 877
rect 2395 843 2433 877
rect 2467 843 2483 877
rect 220 777 254 793
rect 220 709 254 743
rect 220 641 254 667
rect 220 591 254 595
rect 436 777 470 793
rect 436 709 470 743
rect 436 641 470 667
rect 436 591 470 595
rect 546 785 580 793
rect 546 713 580 743
rect 546 641 580 675
rect 546 591 580 607
rect 762 777 796 793
rect 762 709 796 743
rect 762 641 796 643
rect 762 605 796 607
rect 978 785 1012 793
rect 978 713 1012 743
rect 978 641 1012 675
rect 978 591 1012 607
rect 1194 777 1228 793
rect 1194 741 1228 743
rect 1194 641 1228 675
rect 1194 605 1228 607
rect 1304 664 1338 691
rect 1304 589 1338 623
rect 1304 521 1338 553
rect 288 441 303 475
rect 358 441 379 475
rect 427 441 455 475
rect 496 441 531 475
rect 565 441 600 475
rect 641 441 669 475
rect 717 441 738 475
rect 793 441 807 475
rect 869 441 876 475
rect 910 441 911 475
rect 979 441 987 475
rect 1048 441 1063 475
rect 1117 441 1139 475
rect 1186 441 1210 475
rect 1304 453 1338 476
rect 1304 385 1338 399
rect 1304 317 1338 322
rect 1304 279 1338 283
rect 1304 201 1338 215
rect 649 155 687 156
rect 255 121 271 155
rect 315 121 353 155
rect 403 121 467 155
rect 501 121 517 155
rect 577 121 593 155
rect 649 122 683 155
rect 721 122 733 155
rect 627 121 683 122
rect 717 121 733 122
rect 789 121 805 155
rect 856 121 894 155
rect 929 121 945 155
rect 1001 121 1013 155
rect 1051 121 1085 155
rect 1141 121 1157 155
rect 1304 123 1338 147
rect 210 65 244 77
rect 210 -7 244 27
rect 210 -75 244 -41
rect 210 -125 244 -109
rect 316 61 350 77
rect 316 -7 350 27
rect 316 -44 350 -41
rect 316 -116 350 -109
rect 422 65 456 77
rect 422 -7 456 27
rect 422 -75 456 -41
rect 422 -125 456 -109
rect 528 61 562 77
rect 528 -7 562 27
rect 528 -44 562 -41
rect 528 -116 562 -109
rect 638 61 672 77
rect 638 -7 672 -6
rect 638 -44 672 -41
rect 638 -125 672 -109
rect 744 61 778 77
rect 744 -7 778 27
rect 744 -44 778 -41
rect 744 -116 778 -109
rect 850 61 884 77
rect 850 -7 884 27
rect 850 -75 884 -45
rect 850 -125 884 -109
rect 956 61 990 77
rect 956 -7 990 27
rect 956 -44 990 -41
rect 956 -116 990 -109
rect 1062 61 1096 77
rect 1062 -7 1096 27
rect 1062 -75 1096 -45
rect 1062 -125 1096 -109
rect 1168 61 1202 77
rect 1168 -7 1202 27
rect 1168 -44 1202 -41
rect 1168 -116 1202 -109
rect 1304 45 1338 79
rect 1304 -23 1338 11
rect 1304 -91 1338 -57
rect 1304 -159 1338 -125
rect 1304 -209 1338 -193
rect 1520 725 1554 741
rect 1520 657 1554 691
rect 1520 609 1554 623
rect 1520 533 1554 555
rect 1520 457 1554 487
rect 1520 385 1554 419
rect 1520 317 1554 347
rect 1520 249 1554 271
rect 1520 181 1554 194
rect 1520 113 1554 117
rect 1520 74 1554 79
rect 1520 -3 1554 11
rect 1520 -80 1554 -57
rect 1520 -159 1554 -125
rect 1520 -209 1554 -193
rect 1736 664 1770 691
rect 1736 589 1770 623
rect 1736 521 1770 553
rect 1736 453 1770 476
rect 1736 385 1770 399
rect 1736 317 1770 322
rect 1736 279 1770 283
rect 1736 201 1770 215
rect 1736 123 1770 147
rect 1736 45 1770 79
rect 1736 -23 1770 11
rect 1736 -91 1770 -57
rect 1736 -159 1770 -125
rect 1736 -209 1770 -193
rect 1952 725 1986 741
rect 1952 657 1986 691
rect 1952 589 1986 623
rect 1952 521 1986 555
rect 1952 453 1986 487
rect 1952 385 1986 410
rect 1952 317 1986 333
rect 1952 249 1986 256
rect 1952 213 1986 215
rect 1952 136 1986 147
rect 1952 59 1986 79
rect 1952 -19 1986 11
rect 1952 -91 1986 -57
rect 1952 -159 1986 -131
rect 2168 664 2202 691
rect 2168 589 2202 623
rect 2168 521 2202 553
rect 2168 453 2202 476
rect 2168 385 2202 399
rect 2168 317 2202 322
rect 2168 279 2202 283
rect 2168 201 2202 215
rect 2168 123 2202 147
rect 2168 45 2202 79
rect 2168 -23 2202 11
rect 2168 -91 2202 -57
rect 2168 -159 2202 -125
rect 2168 -209 2202 -193
rect 2278 665 2312 691
rect 2278 589 2312 623
rect 2278 521 2312 555
rect 2278 453 2312 479
rect 2278 385 2312 403
rect 2278 317 2312 327
rect 2278 249 2312 251
rect 2278 209 2312 215
rect 2278 133 2312 147
rect 2278 56 2312 79
rect 2278 -21 2312 11
rect 2278 -91 2312 -57
rect 2278 -159 2312 -132
rect 2494 665 2528 691
rect 2494 589 2528 623
rect 2494 521 2528 555
rect 2494 453 2528 479
rect 2494 385 2528 403
rect 2494 317 2528 327
rect 2494 249 2528 251
rect 2494 209 2528 215
rect 2494 133 2528 147
rect 2494 56 2528 79
rect 2494 -21 2528 11
rect 2494 -91 2528 -57
rect 2494 -159 2528 -132
rect 230 -315 246 -281
rect 301 -315 320 -281
rect 372 -315 394 -281
rect 442 -315 468 -281
rect 512 -315 542 -281
rect 582 -315 616 -281
rect 652 -315 688 -281
rect 724 -315 758 -281
rect 798 -315 828 -281
rect 872 -315 898 -281
rect 946 -315 968 -281
rect 1020 -315 1038 -281
rect 1094 -315 1108 -281
rect 1168 -315 1178 -281
rect 1242 -315 1248 -281
rect 1316 -315 1318 -281
rect 1352 -315 1355 -281
rect 1422 -315 1428 -281
rect 1492 -315 1501 -281
rect 1562 -315 1574 -281
rect 1632 -315 1647 -281
rect 1702 -315 1720 -281
rect 1772 -315 1793 -281
rect 1842 -315 1866 -281
rect 1912 -315 1939 -281
rect 1982 -315 2012 -281
rect 2052 -315 2085 -281
rect 2122 -315 2158 -281
rect 2192 -315 2228 -281
rect 2265 -315 2298 -281
rect 2338 -315 2368 -281
rect 2411 -315 2438 -281
rect 2484 -315 2496 -281
<< viali >>
rect 673 3544 677 3578
rect 677 3544 707 3578
rect 750 3544 779 3578
rect 779 3544 784 3578
rect 827 3544 847 3578
rect 847 3544 861 3578
rect 904 3544 915 3578
rect 915 3544 938 3578
rect 981 3544 983 3578
rect 983 3544 1015 3578
rect 1058 3544 1085 3578
rect 1085 3544 1092 3578
rect 1135 3544 1169 3578
rect 1494 3552 1498 3586
rect 1498 3552 1528 3586
rect 1566 3552 1600 3586
rect 1330 3525 1364 3526
rect 1330 3492 1364 3525
rect 674 3446 690 3480
rect 690 3446 708 3480
rect 757 3446 758 3480
rect 758 3446 791 3480
rect 840 3446 860 3480
rect 860 3446 874 3480
rect 922 3446 928 3480
rect 928 3446 956 3480
rect 1004 3446 1030 3480
rect 1030 3446 1038 3480
rect 1086 3446 1098 3480
rect 1098 3446 1120 3480
rect 1168 3446 1200 3480
rect 1200 3446 1202 3480
rect 1694 3514 1728 3534
rect 1694 3500 1728 3514
rect 1330 3435 1364 3454
rect 1414 3446 1430 3480
rect 1430 3446 1448 3480
rect 1486 3446 1498 3480
rect 1498 3446 1520 3480
rect 1694 3446 1728 3462
rect 452 3391 462 3425
rect 462 3391 486 3425
rect 524 3391 530 3425
rect 530 3391 558 3425
rect 1330 3420 1364 3435
rect 1694 3428 1728 3446
rect 1694 3378 1728 3390
rect 746 3340 758 3374
rect 758 3340 780 3374
rect 831 3340 860 3374
rect 860 3340 865 3374
rect 916 3340 928 3374
rect 928 3340 950 3374
rect 1001 3340 1030 3374
rect 1030 3340 1035 3374
rect 1086 3340 1098 3374
rect 1098 3340 1120 3374
rect 1170 3340 1200 3374
rect 1200 3340 1204 3374
rect 1494 3340 1498 3374
rect 1498 3340 1528 3374
rect 1566 3340 1600 3374
rect 1694 3356 1728 3378
rect 1694 3310 1728 3318
rect 1694 3284 1728 3310
rect 666 3230 682 3264
rect 682 3230 700 3264
rect 745 3230 750 3264
rect 750 3230 779 3264
rect 824 3230 852 3264
rect 852 3230 858 3264
rect 903 3230 920 3264
rect 920 3230 937 3264
rect 982 3230 988 3264
rect 988 3230 1016 3264
rect 1061 3230 1090 3264
rect 1090 3230 1095 3264
rect 1140 3230 1158 3264
rect 1158 3230 1174 3264
rect 1219 3230 1226 3264
rect 1226 3230 1253 3264
rect 1297 3230 1328 3264
rect 1328 3230 1331 3264
rect 1375 3230 1396 3264
rect 1396 3230 1409 3264
rect 1453 3230 1464 3264
rect 1464 3230 1487 3264
rect 1694 3242 1728 3246
rect 454 3185 462 3212
rect 462 3185 488 3212
rect 526 3185 530 3212
rect 530 3185 560 3212
rect 1694 3212 1728 3242
rect 454 3178 488 3185
rect 526 3178 560 3185
rect 795 3124 818 3158
rect 818 3124 829 3158
rect 874 3124 886 3158
rect 886 3124 908 3158
rect 953 3124 954 3158
rect 954 3124 987 3158
rect 1032 3124 1056 3158
rect 1056 3124 1066 3158
rect 1111 3124 1124 3158
rect 1124 3124 1145 3158
rect 1190 3124 1192 3158
rect 1192 3124 1224 3158
rect 1269 3124 1294 3158
rect 1294 3124 1303 3158
rect 1348 3124 1362 3158
rect 1362 3124 1382 3158
rect 1426 3124 1430 3158
rect 1430 3124 1460 3158
rect 1504 3124 1532 3158
rect 1532 3124 1538 3158
rect 1582 3124 1600 3158
rect 1600 3124 1616 3158
rect 1694 3140 1728 3174
rect 450 3071 462 3105
rect 462 3071 484 3105
rect 522 3071 530 3105
rect 530 3071 556 3105
rect 1694 3072 1728 3102
rect 1694 3068 1728 3072
rect 666 3018 682 3052
rect 682 3018 700 3052
rect 745 3018 750 3052
rect 750 3018 779 3052
rect 824 3018 852 3052
rect 852 3018 858 3052
rect 903 3018 920 3052
rect 920 3018 937 3052
rect 982 3018 988 3052
rect 988 3018 1016 3052
rect 1061 3018 1090 3052
rect 1090 3018 1095 3052
rect 1140 3018 1158 3052
rect 1158 3018 1174 3052
rect 1219 3018 1226 3052
rect 1226 3018 1253 3052
rect 1297 3018 1328 3052
rect 1328 3018 1331 3052
rect 1375 3018 1396 3052
rect 1396 3018 1409 3052
rect 1453 3018 1464 3052
rect 1464 3018 1487 3052
rect 1694 3004 1728 3029
rect 1694 2995 1728 3004
rect 666 2908 682 2942
rect 682 2908 700 2942
rect 745 2908 750 2942
rect 750 2908 779 2942
rect 824 2908 852 2942
rect 852 2908 858 2942
rect 903 2908 920 2942
rect 920 2908 937 2942
rect 982 2908 988 2942
rect 988 2908 1016 2942
rect 1061 2908 1090 2942
rect 1090 2908 1095 2942
rect 1140 2908 1158 2942
rect 1158 2908 1174 2942
rect 1219 2908 1226 2942
rect 1226 2908 1253 2942
rect 1297 2908 1328 2942
rect 1328 2908 1331 2942
rect 1375 2908 1396 2942
rect 1396 2908 1409 2942
rect 1453 2908 1464 2942
rect 1464 2908 1487 2942
rect 1694 2936 1728 2956
rect 1694 2922 1728 2936
rect 452 2857 462 2891
rect 462 2857 486 2891
rect 524 2857 530 2891
rect 530 2857 558 2891
rect 1694 2868 1728 2883
rect 1694 2849 1728 2868
rect 795 2802 818 2836
rect 818 2802 829 2836
rect 874 2802 886 2836
rect 886 2802 908 2836
rect 953 2802 954 2836
rect 954 2802 987 2836
rect 1032 2802 1056 2836
rect 1056 2802 1066 2836
rect 1111 2802 1124 2836
rect 1124 2802 1145 2836
rect 1190 2802 1192 2836
rect 1192 2802 1224 2836
rect 1269 2802 1294 2836
rect 1294 2802 1303 2836
rect 1348 2802 1362 2836
rect 1362 2802 1382 2836
rect 1426 2802 1430 2836
rect 1430 2802 1460 2836
rect 1504 2802 1532 2836
rect 1532 2802 1538 2836
rect 1582 2802 1600 2836
rect 1600 2802 1616 2836
rect 1694 2800 1728 2810
rect 530 2741 564 2765
rect 530 2731 564 2741
rect 1694 2776 1728 2800
rect 1694 2732 1728 2737
rect 666 2696 682 2730
rect 682 2696 700 2730
rect 745 2696 750 2730
rect 750 2696 779 2730
rect 824 2696 852 2730
rect 852 2696 858 2730
rect 903 2696 920 2730
rect 920 2696 937 2730
rect 982 2696 988 2730
rect 988 2696 1016 2730
rect 1061 2696 1090 2730
rect 1090 2696 1095 2730
rect 1140 2696 1158 2730
rect 1158 2696 1174 2730
rect 1219 2696 1226 2730
rect 1226 2696 1253 2730
rect 1297 2696 1328 2730
rect 1328 2696 1331 2730
rect 1375 2696 1396 2730
rect 1396 2696 1409 2730
rect 1453 2696 1464 2730
rect 1464 2696 1487 2730
rect 1694 2703 1728 2732
rect 530 2677 564 2683
rect 530 2649 564 2677
rect 1694 2630 1728 2664
rect 530 2579 564 2601
rect 795 2590 818 2624
rect 818 2590 829 2624
rect 874 2590 886 2624
rect 886 2590 908 2624
rect 953 2590 954 2624
rect 954 2590 987 2624
rect 1032 2590 1056 2624
rect 1056 2590 1066 2624
rect 1111 2590 1124 2624
rect 1124 2590 1145 2624
rect 1190 2590 1192 2624
rect 1192 2590 1224 2624
rect 1269 2590 1294 2624
rect 1294 2590 1303 2624
rect 1348 2590 1362 2624
rect 1362 2590 1382 2624
rect 1426 2590 1430 2624
rect 1430 2590 1460 2624
rect 1504 2590 1532 2624
rect 1532 2590 1538 2624
rect 1582 2590 1600 2624
rect 1600 2590 1616 2624
rect 530 2567 564 2579
rect 666 2484 682 2518
rect 682 2484 700 2518
rect 745 2484 750 2518
rect 750 2484 779 2518
rect 824 2484 852 2518
rect 852 2484 858 2518
rect 903 2484 920 2518
rect 920 2484 937 2518
rect 982 2484 988 2518
rect 988 2484 1016 2518
rect 1061 2484 1090 2518
rect 1090 2484 1095 2518
rect 1140 2484 1158 2518
rect 1158 2484 1174 2518
rect 1219 2484 1226 2518
rect 1226 2484 1253 2518
rect 1297 2484 1328 2518
rect 1328 2484 1331 2518
rect 1375 2484 1396 2518
rect 1396 2484 1409 2518
rect 1453 2484 1464 2518
rect 1464 2484 1487 2518
rect 699 1968 722 2002
rect 722 1968 733 2002
rect 776 1968 790 2002
rect 790 1968 810 2002
rect 853 1968 858 2002
rect 858 1968 887 2002
rect 930 1968 960 2002
rect 960 1968 964 2002
rect 1007 1968 1028 2002
rect 1028 1968 1041 2002
rect 1084 1968 1096 2002
rect 1096 1968 1118 2002
rect 1161 1968 1164 2002
rect 1164 1968 1195 2002
rect 1238 1968 1266 2002
rect 1266 1968 1272 2002
rect 1314 1968 1334 2002
rect 1334 1968 1348 2002
rect 1390 1968 1402 2002
rect 1402 1968 1424 2002
rect 1466 1968 1470 2002
rect 1470 1968 1500 2002
rect 1542 1968 1572 2002
rect 1572 1968 1576 2002
rect 1716 1963 1750 1997
rect 560 1907 594 1915
rect 560 1881 594 1907
rect 560 1789 594 1823
rect 1716 1903 1750 1925
rect 1716 1891 1750 1903
rect 1716 1835 1750 1853
rect 1716 1819 1750 1835
rect 699 1752 722 1786
rect 722 1752 733 1786
rect 777 1752 790 1786
rect 790 1752 811 1786
rect 855 1752 858 1786
rect 858 1752 889 1786
rect 933 1752 960 1786
rect 960 1752 967 1786
rect 1011 1752 1028 1786
rect 1028 1752 1045 1786
rect 1089 1752 1096 1786
rect 1096 1752 1123 1786
rect 1167 1752 1198 1786
rect 1198 1752 1201 1786
rect 1245 1752 1266 1786
rect 1266 1752 1279 1786
rect 1322 1752 1334 1786
rect 1334 1752 1356 1786
rect 1399 1752 1402 1786
rect 1402 1752 1433 1786
rect 1476 1752 1504 1786
rect 1504 1752 1510 1786
rect 1553 1752 1572 1786
rect 1572 1752 1587 1786
rect 1716 1767 1750 1781
rect 560 1709 594 1731
rect 560 1697 594 1709
rect 560 1631 594 1638
rect 560 1604 594 1631
rect 1716 1747 1750 1767
rect 1716 1699 1750 1709
rect 1716 1675 1750 1699
rect 1716 1631 1750 1636
rect 1716 1602 1750 1631
rect 699 1536 722 1570
rect 722 1536 733 1570
rect 777 1536 790 1570
rect 790 1536 811 1570
rect 855 1536 858 1570
rect 858 1536 889 1570
rect 933 1536 960 1570
rect 960 1536 967 1570
rect 1011 1536 1028 1570
rect 1028 1536 1045 1570
rect 1089 1536 1096 1570
rect 1096 1536 1123 1570
rect 1167 1536 1198 1570
rect 1198 1536 1201 1570
rect 1245 1536 1266 1570
rect 1266 1536 1279 1570
rect 1322 1536 1334 1570
rect 1334 1536 1356 1570
rect 1399 1536 1402 1570
rect 1402 1536 1433 1570
rect 1476 1536 1504 1570
rect 1504 1536 1510 1570
rect 1553 1536 1572 1570
rect 1572 1536 1587 1570
rect 1716 1529 1750 1563
rect 291 843 315 877
rect 315 843 325 877
rect 363 843 375 877
rect 375 843 397 877
rect 631 843 641 877
rect 641 843 665 877
rect 711 843 717 877
rect 717 843 745 877
rect 791 843 792 877
rect 792 843 825 877
rect 871 843 905 877
rect 950 843 983 877
rect 983 843 984 877
rect 1029 843 1058 877
rect 1058 843 1063 877
rect 1108 843 1133 877
rect 1133 843 1142 877
rect 1369 843 1399 877
rect 1399 843 1403 877
rect 1444 843 1474 877
rect 1474 843 1478 877
rect 1519 843 1549 877
rect 1549 843 1553 877
rect 1594 843 1623 877
rect 1623 843 1628 877
rect 1668 843 1697 877
rect 1697 843 1702 877
rect 1742 843 1771 877
rect 1771 843 1776 877
rect 1816 843 1845 877
rect 1845 843 1850 877
rect 1890 843 1919 877
rect 1919 843 1924 877
rect 1964 843 1993 877
rect 1993 843 1998 877
rect 2038 843 2067 877
rect 2067 843 2072 877
rect 2112 843 2141 877
rect 2141 843 2146 877
rect 2361 843 2373 877
rect 2373 843 2395 877
rect 2433 843 2467 877
rect 220 675 254 701
rect 220 667 254 675
rect 220 607 254 629
rect 220 595 254 607
rect 436 675 470 701
rect 436 667 470 675
rect 436 607 470 629
rect 436 595 470 607
rect 546 777 580 785
rect 546 751 580 777
rect 546 709 580 713
rect 546 679 580 709
rect 762 675 796 677
rect 762 643 796 675
rect 762 571 796 605
rect 978 777 1012 785
rect 978 751 1012 777
rect 978 709 1012 713
rect 978 679 1012 709
rect 1194 709 1228 741
rect 1194 707 1228 709
rect 1194 571 1228 605
rect 1304 725 1338 741
rect 1304 707 1338 725
rect 1304 657 1338 664
rect 1304 630 1338 657
rect 1304 555 1338 587
rect 1304 553 1338 555
rect 1304 487 1338 510
rect 1304 476 1338 487
rect 226 441 254 475
rect 254 441 260 475
rect 303 441 324 475
rect 324 441 337 475
rect 379 441 393 475
rect 393 441 413 475
rect 455 441 462 475
rect 462 441 489 475
rect 531 441 565 475
rect 607 441 634 475
rect 634 441 641 475
rect 683 441 703 475
rect 703 441 717 475
rect 759 441 772 475
rect 772 441 793 475
rect 835 441 841 475
rect 841 441 869 475
rect 911 441 945 475
rect 987 441 1014 475
rect 1014 441 1021 475
rect 1063 441 1083 475
rect 1083 441 1097 475
rect 1139 441 1152 475
rect 1152 441 1173 475
rect 1304 419 1338 433
rect 1304 399 1338 419
rect 1304 351 1338 356
rect 1304 322 1338 351
rect 1304 249 1338 279
rect 1304 245 1338 249
rect 1304 181 1338 201
rect 1304 167 1338 181
rect 615 155 649 156
rect 687 155 721 156
rect 281 121 305 155
rect 305 121 315 155
rect 353 121 369 155
rect 369 121 387 155
rect 615 122 627 155
rect 627 122 649 155
rect 687 122 717 155
rect 717 122 721 155
rect 822 121 839 155
rect 839 121 856 155
rect 894 121 895 155
rect 895 121 928 155
rect 1013 121 1017 155
rect 1017 121 1047 155
rect 1085 121 1107 155
rect 1107 121 1119 155
rect 1304 113 1338 123
rect 1304 89 1338 113
rect 210 61 244 65
rect 210 31 244 61
rect 210 -41 244 -7
rect 316 -75 350 -44
rect 316 -78 350 -75
rect 316 -150 350 -116
rect 422 61 456 65
rect 422 31 456 61
rect 422 -41 456 -7
rect 528 -75 562 -44
rect 528 -78 562 -75
rect 528 -150 562 -116
rect 638 27 672 28
rect 638 -6 672 27
rect 638 -75 672 -44
rect 638 -78 672 -75
rect 744 -75 778 -44
rect 744 -78 778 -75
rect 744 -150 778 -116
rect 850 27 884 61
rect 850 -41 884 -11
rect 850 -45 884 -41
rect 956 -75 990 -44
rect 956 -78 990 -75
rect 956 -150 990 -116
rect 1062 27 1096 61
rect 1062 -41 1096 -11
rect 1062 -45 1096 -41
rect 1168 -75 1202 -44
rect 1168 -78 1202 -75
rect 1168 -150 1202 -116
rect 1304 11 1338 45
rect 1520 589 1554 609
rect 1520 575 1554 589
rect 1520 521 1554 533
rect 1520 499 1554 521
rect 1520 453 1554 457
rect 1520 423 1554 453
rect 1520 351 1554 381
rect 1520 347 1554 351
rect 1520 283 1554 305
rect 1520 271 1554 283
rect 1520 215 1554 228
rect 1520 194 1554 215
rect 1520 147 1554 151
rect 1520 117 1554 147
rect 1520 45 1554 74
rect 1520 40 1554 45
rect 1520 -23 1554 -3
rect 1520 -37 1554 -23
rect 1520 -91 1554 -80
rect 1520 -114 1554 -91
rect 1736 725 1770 741
rect 1736 707 1770 725
rect 1736 657 1770 664
rect 1736 630 1770 657
rect 1736 555 1770 587
rect 1736 553 1770 555
rect 1736 487 1770 510
rect 1736 476 1770 487
rect 1736 419 1770 433
rect 1736 399 1770 419
rect 1736 351 1770 356
rect 1736 322 1770 351
rect 1736 249 1770 279
rect 1736 245 1770 249
rect 1736 181 1770 201
rect 1736 167 1770 181
rect 1736 113 1770 123
rect 1736 89 1770 113
rect 1736 11 1770 45
rect 1952 487 1986 521
rect 1952 419 1986 444
rect 1952 410 1986 419
rect 1952 351 1986 367
rect 1952 333 1986 351
rect 1952 283 1986 290
rect 1952 256 1986 283
rect 1952 181 1986 213
rect 1952 179 1986 181
rect 1952 113 1986 136
rect 1952 102 1986 113
rect 1952 45 1986 59
rect 1952 25 1986 45
rect 1952 -23 1986 -19
rect 1952 -53 1986 -23
rect 1952 -125 1986 -97
rect 1952 -131 1986 -125
rect 1952 -193 1986 -175
rect 1952 -209 1986 -193
rect 2168 725 2202 741
rect 2168 707 2202 725
rect 2168 657 2202 664
rect 2168 630 2202 657
rect 2168 555 2202 587
rect 2168 553 2202 555
rect 2168 487 2202 510
rect 2168 476 2202 487
rect 2168 419 2202 433
rect 2168 399 2202 419
rect 2168 351 2202 356
rect 2168 322 2202 351
rect 2168 249 2202 279
rect 2168 245 2202 249
rect 2168 181 2202 201
rect 2168 167 2202 181
rect 2168 113 2202 123
rect 2168 89 2202 113
rect 2168 11 2202 45
rect 2278 725 2312 741
rect 2278 707 2312 725
rect 2278 657 2312 665
rect 2278 631 2312 657
rect 2278 555 2312 589
rect 2278 487 2312 513
rect 2278 479 2312 487
rect 2278 419 2312 437
rect 2278 403 2312 419
rect 2278 351 2312 361
rect 2278 327 2312 351
rect 2278 283 2312 285
rect 2278 251 2312 283
rect 2278 181 2312 209
rect 2278 175 2312 181
rect 2278 113 2312 133
rect 2278 99 2312 113
rect 2278 45 2312 56
rect 2278 22 2312 45
rect 2278 -23 2312 -21
rect 2278 -55 2312 -23
rect 2278 -125 2312 -98
rect 2278 -132 2312 -125
rect 2278 -193 2312 -175
rect 2278 -209 2312 -193
rect 2494 725 2528 741
rect 2494 707 2528 725
rect 2494 657 2528 665
rect 2494 631 2528 657
rect 2494 555 2528 589
rect 2494 487 2528 513
rect 2494 479 2528 487
rect 2494 419 2528 437
rect 2494 403 2528 419
rect 2494 351 2528 361
rect 2494 327 2528 351
rect 2494 283 2528 285
rect 2494 251 2528 283
rect 2494 181 2528 209
rect 2494 175 2528 181
rect 2494 113 2528 133
rect 2494 99 2528 113
rect 2494 45 2528 56
rect 2494 22 2528 45
rect 2494 -23 2528 -21
rect 2494 -55 2528 -23
rect 2494 -125 2528 -98
rect 2494 -132 2528 -125
rect 2494 -193 2528 -175
rect 2494 -209 2528 -193
rect 172 -315 196 -281
rect 196 -315 206 -281
rect 246 -315 267 -281
rect 267 -315 280 -281
rect 320 -315 338 -281
rect 338 -315 354 -281
rect 394 -315 408 -281
rect 408 -315 428 -281
rect 468 -315 478 -281
rect 478 -315 502 -281
rect 542 -315 548 -281
rect 548 -315 576 -281
rect 616 -315 618 -281
rect 618 -315 650 -281
rect 690 -315 722 -281
rect 722 -315 724 -281
rect 764 -315 792 -281
rect 792 -315 798 -281
rect 838 -315 862 -281
rect 862 -315 872 -281
rect 912 -315 932 -281
rect 932 -315 946 -281
rect 986 -315 1002 -281
rect 1002 -315 1020 -281
rect 1060 -315 1072 -281
rect 1072 -315 1094 -281
rect 1134 -315 1142 -281
rect 1142 -315 1168 -281
rect 1208 -315 1212 -281
rect 1212 -315 1242 -281
rect 1282 -315 1316 -281
rect 1355 -315 1388 -281
rect 1388 -315 1389 -281
rect 1428 -315 1458 -281
rect 1458 -315 1462 -281
rect 1501 -315 1528 -281
rect 1528 -315 1535 -281
rect 1574 -315 1598 -281
rect 1598 -315 1608 -281
rect 1647 -315 1668 -281
rect 1668 -315 1681 -281
rect 1720 -315 1738 -281
rect 1738 -315 1754 -281
rect 1793 -315 1808 -281
rect 1808 -315 1827 -281
rect 1866 -315 1878 -281
rect 1878 -315 1900 -281
rect 1939 -315 1948 -281
rect 1948 -315 1973 -281
rect 2012 -315 2018 -281
rect 2018 -315 2046 -281
rect 2085 -315 2088 -281
rect 2088 -315 2119 -281
rect 2158 -315 2192 -281
rect 2231 -315 2262 -281
rect 2262 -315 2265 -281
rect 2304 -315 2332 -281
rect 2332 -315 2338 -281
rect 2377 -315 2402 -281
rect 2402 -315 2411 -281
rect 2450 -315 2472 -281
rect 2472 -315 2484 -281
<< metal1 >>
rect 1683 3639 1799 3645
rect 1482 3586 1612 3592
rect 661 3578 1214 3584
rect 661 3577 673 3578
rect 707 3577 750 3578
rect 784 3577 827 3578
rect 661 3525 671 3577
rect 723 3544 750 3577
rect 820 3544 827 3577
rect 861 3577 904 3578
rect 938 3577 981 3578
rect 861 3544 865 3577
rect 938 3544 962 3577
rect 1015 3544 1058 3578
rect 1092 3577 1135 3578
rect 1169 3577 1214 3578
rect 1111 3544 1135 3577
rect 723 3525 768 3544
rect 820 3525 865 3544
rect 917 3525 962 3544
rect 1014 3525 1059 3544
rect 1111 3525 1156 3544
rect 1208 3525 1214 3577
rect 1482 3552 1494 3586
rect 1528 3552 1566 3586
rect 1600 3552 1612 3586
rect 1482 3546 1612 3552
tri 1529 3538 1537 3546 ne
rect 1537 3538 1612 3546
rect 661 3480 1214 3525
rect 1324 3526 1370 3538
tri 1537 3534 1541 3538 ne
rect 1541 3534 1612 3538
tri 1322 3492 1324 3494 se
rect 1324 3492 1330 3526
rect 1364 3492 1370 3526
tri 1541 3517 1558 3534 ne
rect 1558 3517 1612 3534
tri 1558 3512 1563 3517 ne
tri 1316 3486 1322 3492 se
rect 1322 3486 1370 3492
tri 1310 3480 1316 3486 se
rect 1316 3480 1370 3486
rect 661 3446 674 3480
rect 708 3446 757 3480
rect 791 3446 840 3480
rect 874 3446 922 3480
rect 956 3446 1004 3480
rect 1038 3446 1086 3480
rect 1120 3446 1168 3480
rect 1202 3446 1214 3480
tri 1290 3460 1310 3480 se
rect 1310 3460 1370 3480
rect 661 3440 1214 3446
rect 440 3382 448 3434
rect 500 3382 512 3434
rect 564 3382 570 3434
rect 1242 3408 1248 3460
rect 1300 3408 1312 3460
rect 1364 3408 1370 3460
rect 1402 3436 1410 3488
rect 1462 3436 1474 3488
rect 1526 3436 1532 3488
tri 1557 3408 1563 3414 se
rect 1563 3408 1612 3517
tri 1539 3390 1557 3408 se
rect 1557 3390 1612 3408
tri 1531 3382 1539 3390 se
rect 1539 3382 1612 3390
tri 1529 3380 1531 3382 se
rect 1531 3380 1612 3382
rect 734 3374 1612 3380
rect 734 3340 746 3374
rect 780 3340 831 3374
rect 865 3340 916 3374
rect 950 3340 1001 3374
rect 1035 3340 1086 3374
rect 1120 3340 1170 3374
rect 1204 3340 1494 3374
rect 1528 3340 1566 3374
rect 1600 3340 1612 3374
rect 734 3334 1612 3340
rect 1683 3500 1694 3523
rect 1728 3500 1799 3523
rect 1683 3462 1799 3500
rect 1683 3428 1694 3462
rect 1728 3428 1799 3462
rect 1683 3412 1799 3428
rect 1683 3390 1707 3412
rect 1683 3356 1694 3390
rect 1759 3360 1799 3412
rect 1728 3356 1799 3360
rect 1683 3329 1799 3356
rect 1683 3318 1707 3329
rect 1683 3284 1694 3318
rect 1683 3277 1707 3284
rect 1759 3277 1799 3329
rect 654 3264 1032 3273
rect 1084 3264 1096 3273
rect 1148 3264 1499 3273
rect 654 3230 666 3264
rect 700 3230 745 3264
rect 779 3230 824 3264
rect 858 3230 903 3264
rect 937 3230 982 3264
rect 1016 3230 1032 3264
rect 1095 3230 1096 3264
rect 1174 3230 1219 3264
rect 1253 3230 1297 3264
rect 1331 3230 1375 3264
rect 1409 3230 1453 3264
rect 1487 3230 1499 3264
rect 654 3221 1032 3230
rect 1084 3221 1096 3230
rect 1148 3221 1499 3230
rect 1683 3246 1799 3277
rect 442 3212 615 3218
tri 615 3212 621 3218 sw
rect 1683 3212 1694 3246
rect 442 3178 454 3212
rect 488 3178 526 3212
rect 560 3178 621 3212
rect 442 3174 621 3178
tri 621 3174 659 3212 sw
tri 1659 3174 1683 3198 se
rect 1683 3194 1707 3212
rect 1759 3194 1799 3246
rect 1683 3174 1799 3194
rect 442 3172 659 3174
tri 595 3161 606 3172 ne
rect 606 3164 659 3172
tri 659 3164 669 3174 sw
tri 1649 3164 1659 3174 se
rect 1659 3164 1694 3174
rect 606 3161 669 3164
tri 669 3161 672 3164 sw
tri 606 3158 609 3161 ne
rect 609 3158 672 3161
tri 609 3152 615 3158 ne
rect 615 3152 672 3158
tri 615 3141 626 3152 ne
rect 438 3062 444 3114
rect 496 3062 508 3114
rect 560 3062 568 3114
rect 626 3068 672 3152
rect 783 3158 1694 3164
rect 1728 3163 1799 3174
rect 783 3124 795 3158
rect 829 3124 874 3158
rect 908 3124 953 3158
rect 987 3124 1032 3158
rect 1066 3124 1111 3158
rect 1145 3124 1190 3158
rect 1224 3124 1269 3158
rect 1303 3124 1348 3158
rect 1382 3124 1426 3158
rect 1460 3124 1504 3158
rect 1538 3124 1582 3158
rect 1616 3140 1694 3158
rect 1616 3124 1707 3140
rect 783 3118 1707 3124
tri 1539 3102 1555 3118 ne
rect 1555 3111 1707 3118
rect 1759 3111 1799 3163
rect 1555 3102 1799 3111
tri 1555 3095 1562 3102 ne
rect 1562 3095 1694 3102
tri 672 3068 699 3095 sw
tri 1562 3084 1573 3095 ne
rect 1573 3068 1694 3095
rect 1728 3080 1799 3102
rect 626 3062 699 3068
tri 699 3062 705 3068 sw
rect 626 3061 705 3062
tri 705 3061 706 3062 sw
rect 626 3052 876 3061
rect 928 3052 940 3061
rect 992 3052 1499 3061
rect 626 3018 666 3052
rect 700 3018 745 3052
rect 779 3018 824 3052
rect 858 3018 876 3052
rect 937 3018 940 3052
rect 1016 3018 1061 3052
rect 1095 3018 1140 3052
rect 1174 3018 1219 3052
rect 1253 3018 1297 3052
rect 1331 3018 1375 3052
rect 1409 3018 1453 3052
rect 1487 3018 1499 3052
rect 626 3009 876 3018
rect 928 3009 940 3018
rect 992 3009 1499 3018
rect 1573 3029 1707 3068
rect 1573 2995 1694 3029
rect 1759 3028 1799 3080
rect 1728 2997 1799 3028
rect 1573 2956 1707 2995
rect 654 2942 708 2951
rect 760 2942 772 2951
rect 824 2942 1499 2951
rect 654 2908 666 2942
rect 700 2908 708 2942
rect 858 2908 903 2942
rect 937 2908 982 2942
rect 1016 2908 1061 2942
rect 1095 2908 1140 2942
rect 1174 2908 1219 2942
rect 1253 2908 1297 2942
rect 1331 2908 1375 2942
rect 1409 2908 1453 2942
rect 1487 2908 1499 2942
rect 654 2899 708 2908
rect 760 2899 772 2908
rect 824 2899 1499 2908
rect 1573 2922 1694 2956
rect 1759 2945 1799 2997
rect 1728 2922 1799 2945
rect 1573 2914 1799 2922
rect 440 2847 448 2899
rect 500 2847 512 2899
rect 564 2847 573 2899
rect 1573 2883 1707 2914
tri 1546 2849 1573 2876 se
rect 1573 2849 1694 2883
rect 1759 2862 1799 2914
rect 1728 2849 1799 2862
tri 487 2842 492 2847 ne
rect 492 2842 573 2847
tri 1539 2842 1546 2849 se
rect 1546 2842 1799 2849
tri 492 2836 498 2842 ne
rect 498 2836 573 2842
tri 498 2813 521 2836 ne
rect 521 2765 573 2836
rect 783 2836 1799 2842
rect 783 2802 795 2836
rect 829 2802 874 2836
rect 908 2802 953 2836
rect 987 2802 1032 2836
rect 1066 2802 1111 2836
rect 1145 2802 1190 2836
rect 1224 2802 1269 2836
rect 1303 2802 1348 2836
rect 1382 2802 1426 2836
rect 1460 2802 1504 2836
rect 1538 2802 1582 2836
rect 1616 2831 1799 2836
rect 1616 2810 1707 2831
rect 1616 2802 1694 2810
rect 783 2796 1694 2802
tri 1539 2776 1559 2796 ne
rect 1559 2776 1694 2796
rect 1759 2779 1799 2831
rect 1728 2776 1799 2779
rect 521 2731 530 2765
rect 564 2731 573 2765
tri 1559 2762 1573 2776 ne
rect 1573 2748 1799 2776
rect 521 2683 573 2731
rect 521 2677 530 2683
rect 564 2677 573 2683
rect 521 2613 573 2625
rect 521 2555 573 2561
rect 654 2730 1180 2739
rect 1232 2730 1244 2739
rect 1296 2730 1499 2739
rect 654 2696 666 2730
rect 700 2696 745 2730
rect 779 2696 824 2730
rect 858 2696 903 2730
rect 937 2696 982 2730
rect 1016 2696 1061 2730
rect 1095 2696 1140 2730
rect 1174 2696 1180 2730
rect 1296 2696 1297 2730
rect 1331 2696 1375 2730
rect 1409 2696 1453 2730
rect 1487 2696 1499 2730
rect 654 2687 1180 2696
rect 1232 2687 1244 2696
rect 1296 2687 1499 2696
rect 1573 2737 1707 2748
rect 1573 2703 1694 2737
rect 1573 2696 1707 2703
rect 1759 2696 1799 2748
rect 654 2664 743 2687
tri 743 2664 766 2687 nw
rect 1573 2665 1799 2696
rect 1573 2664 1707 2665
rect 654 2555 732 2664
tri 732 2653 743 2664 nw
tri 1562 2653 1573 2664 se
rect 1573 2653 1694 2664
tri 1539 2630 1562 2653 se
rect 1562 2630 1694 2653
rect 783 2624 1707 2630
rect 783 2590 795 2624
rect 829 2590 874 2624
rect 908 2590 953 2624
rect 987 2590 1032 2624
rect 1066 2590 1111 2624
rect 1145 2590 1190 2624
rect 1224 2590 1269 2624
rect 1303 2590 1348 2624
rect 1382 2590 1426 2624
rect 1460 2590 1504 2624
rect 1538 2590 1582 2624
rect 1616 2613 1707 2624
rect 1759 2613 1799 2665
rect 1616 2590 1799 2613
rect 783 2584 1799 2590
tri 1539 2561 1562 2584 ne
rect 1562 2582 1799 2584
rect 1562 2561 1707 2582
tri 732 2555 738 2561 sw
tri 1562 2555 1568 2561 ne
rect 1568 2555 1707 2561
rect 654 2527 738 2555
tri 738 2527 766 2555 sw
tri 1568 2550 1573 2555 ne
rect 1573 2530 1707 2555
rect 1759 2530 1799 2582
rect 654 2518 1180 2527
rect 1232 2518 1244 2527
rect 1296 2518 1499 2527
rect 654 2484 666 2518
rect 700 2484 745 2518
rect 779 2484 824 2518
rect 858 2484 903 2518
rect 937 2484 982 2518
rect 1016 2484 1061 2518
rect 1095 2484 1140 2518
rect 1174 2484 1180 2518
rect 1296 2484 1297 2518
rect 1331 2484 1375 2518
rect 1409 2484 1453 2518
rect 1487 2484 1499 2518
rect 654 2475 1180 2484
rect 1232 2475 1244 2484
rect 1296 2475 1499 2484
rect 1573 2498 1799 2530
rect 1573 2446 1707 2498
rect 1759 2446 1799 2498
rect 1573 2440 1799 2446
rect 478 2266 527 2318
rect 579 2266 591 2318
rect 643 2266 788 2318
rect 840 2266 852 2318
rect 904 2266 1636 2318
rect 474 2182 480 2234
rect 532 2182 544 2234
rect 596 2182 1822 2234
rect 1874 2182 1886 2234
rect 1938 2182 1944 2234
rect 687 2002 1180 2011
rect 1232 2002 1244 2011
rect 1296 2002 1588 2011
rect 687 1968 699 2002
rect 733 1968 776 2002
rect 810 1968 853 2002
rect 887 1968 930 2002
rect 964 1968 1007 2002
rect 1041 1968 1084 2002
rect 1118 1968 1161 2002
rect 1232 1968 1238 2002
rect 1296 1968 1314 2002
rect 1348 1968 1390 2002
rect 1424 1968 1466 2002
rect 1500 1968 1542 2002
rect 1576 1968 1588 2002
rect 687 1959 1180 1968
rect 1232 1959 1244 1968
rect 1296 1959 1588 1968
rect 1707 2003 1759 2009
rect 1707 1937 1759 1951
rect 550 1921 602 1927
rect 550 1857 602 1869
rect 1330 1868 1382 1874
rect 866 1843 918 1849
tri 857 1819 866 1828 se
rect 550 1789 560 1805
rect 594 1789 602 1805
tri 832 1794 857 1819 se
rect 857 1794 866 1819
rect 550 1731 602 1789
rect 687 1791 866 1794
tri 918 1819 927 1828 sw
tri 1321 1819 1330 1828 se
rect 918 1794 927 1819
tri 927 1794 952 1819 sw
tri 1296 1794 1321 1819 se
rect 1321 1816 1330 1819
rect 1707 1871 1759 1885
tri 1382 1819 1391 1828 sw
rect 1382 1816 1391 1819
rect 1321 1804 1391 1816
rect 1321 1794 1330 1804
rect 918 1791 1330 1794
rect 687 1786 1330 1791
rect 1382 1794 1391 1804
tri 1391 1794 1416 1819 sw
rect 1707 1805 1759 1819
rect 1382 1786 1496 1794
rect 1548 1786 1560 1794
rect 687 1752 699 1786
rect 733 1752 777 1786
rect 811 1752 855 1786
rect 889 1779 933 1786
rect 918 1752 933 1779
rect 967 1752 1011 1786
rect 1045 1752 1089 1786
rect 1123 1752 1167 1786
rect 1201 1752 1245 1786
rect 1279 1752 1322 1786
rect 1382 1752 1399 1786
rect 1433 1752 1476 1786
rect 1548 1752 1553 1786
rect 687 1742 866 1752
rect 550 1697 560 1731
rect 594 1697 602 1731
tri 845 1721 866 1742 ne
rect 918 1742 1496 1752
rect 1548 1742 1560 1752
rect 1612 1742 1618 1794
rect 1707 1747 1716 1753
rect 1750 1747 1759 1753
rect 866 1721 918 1727
tri 918 1721 939 1742 nw
rect 1707 1739 1759 1747
rect 550 1638 602 1697
rect 550 1604 560 1638
rect 594 1604 602 1638
rect 550 1592 602 1604
rect 1707 1675 1716 1687
rect 1750 1675 1759 1687
rect 1707 1672 1759 1675
rect 1707 1605 1716 1620
rect 1750 1605 1759 1620
rect 687 1570 1180 1579
rect 687 1536 699 1570
rect 733 1536 777 1570
rect 811 1536 855 1570
rect 889 1536 933 1570
rect 967 1536 1011 1570
rect 1045 1536 1089 1570
rect 1123 1536 1167 1570
rect 687 1527 1180 1536
rect 1232 1527 1244 1579
rect 1296 1570 1599 1579
rect 1296 1536 1322 1570
rect 1356 1536 1399 1570
rect 1433 1536 1476 1570
rect 1510 1536 1553 1570
rect 1587 1536 1599 1570
rect 1296 1527 1599 1536
rect 1707 1529 1716 1553
rect 1750 1529 1759 1553
rect 341 1520 393 1526
rect 1707 1517 1759 1529
rect 341 1456 393 1468
tri 393 1450 427 1484 sw
rect 393 1404 533 1450
rect 341 1398 533 1404
rect 585 1398 597 1450
rect 649 1398 1340 1450
rect 1392 1398 1404 1450
rect 1456 1398 1462 1450
rect 421 1318 427 1370
rect 479 1318 491 1370
rect 543 1318 952 1370
rect 1004 1318 1016 1370
rect 1068 1318 1074 1370
rect 204 1238 210 1290
rect 262 1238 274 1290
rect 326 1238 1108 1290
rect 1160 1238 1172 1290
rect 1224 1238 1944 1290
rect 782 1090 788 1142
rect 840 1090 852 1142
rect 904 1090 1109 1142
rect 1161 1090 1173 1142
rect 1225 1090 1231 1142
rect 279 877 476 883
rect 279 843 291 877
rect 325 843 363 877
rect 397 843 476 877
rect 279 837 476 843
tri 396 803 430 837 ne
rect 214 701 260 713
rect 214 667 220 701
rect 254 667 260 701
rect 214 630 260 667
rect 430 701 476 837
rect 619 877 872 886
rect 619 843 631 877
rect 665 843 711 877
rect 745 843 791 877
rect 825 843 871 877
rect 619 834 872 843
rect 924 834 936 886
rect 988 877 1154 886
rect 988 843 1029 877
rect 1063 843 1108 877
rect 1142 843 1154 877
rect 988 834 1154 843
rect 1357 877 1822 886
rect 1357 843 1369 877
rect 1403 843 1444 877
rect 1478 843 1519 877
rect 1553 843 1594 877
rect 1628 843 1668 877
rect 1702 843 1742 877
rect 1776 843 1816 877
rect 1357 834 1822 843
rect 1874 834 1886 886
rect 1938 877 2158 886
rect 1938 843 1964 877
rect 1998 843 2038 877
rect 2072 843 2112 877
rect 2146 843 2158 877
rect 1938 834 2158 843
rect 2349 877 2534 883
rect 2349 843 2361 877
rect 2395 843 2433 877
rect 2467 843 2534 877
rect 2349 837 2534 843
tri 2454 834 2457 837 ne
rect 2457 834 2534 837
tri 2457 803 2488 834 ne
rect 430 667 436 701
rect 470 667 476 701
rect 540 785 1018 797
rect 540 751 546 785
rect 580 784 978 785
rect 580 751 708 784
rect 540 732 708 751
rect 760 732 772 784
rect 824 751 978 784
rect 1012 751 1018 785
rect 824 732 1018 751
rect 540 721 1018 732
rect 540 713 612 721
tri 612 713 620 721 nw
tri 938 713 946 721 ne
rect 946 713 1018 721
rect 540 679 546 713
rect 580 691 590 713
tri 590 691 612 713 nw
tri 946 691 968 713 ne
rect 968 691 978 713
rect 580 689 588 691
tri 588 689 590 691 nw
tri 968 689 970 691 ne
rect 970 689 978 691
rect 580 679 586 689
tri 586 687 588 689 nw
rect 540 667 586 679
rect 756 677 802 689
tri 970 687 972 689 ne
tri 260 630 264 634 sw
tri 426 630 430 634 se
rect 430 630 476 667
rect 214 629 264 630
tri 264 629 265 630 sw
tri 425 629 426 630 se
rect 426 629 476 630
rect 214 595 220 629
rect 254 600 265 629
tri 265 600 294 629 sw
tri 396 600 425 629 se
rect 425 600 436 629
rect 254 595 436 600
rect 470 595 476 629
rect 214 510 476 595
rect 756 643 762 677
rect 796 667 802 677
rect 972 679 978 689
rect 1012 679 1018 713
tri 802 667 808 673 sw
rect 972 667 1018 679
rect 1188 741 2208 753
rect 1188 707 1194 741
rect 1228 707 1304 741
rect 1338 707 1736 741
rect 1770 707 2168 741
rect 2202 707 2208 741
tri 1182 667 1188 673 se
rect 1188 667 2208 707
rect 796 665 808 667
tri 808 665 810 667 sw
tri 1180 665 1182 667 se
rect 1182 665 2208 667
rect 796 664 810 665
tri 810 664 811 665 sw
tri 1179 664 1180 665 se
rect 1180 664 2208 665
rect 796 643 811 664
rect 756 639 811 643
tri 811 639 836 664 sw
tri 1154 639 1179 664 se
rect 1179 639 1304 664
rect 756 630 1304 639
rect 1338 653 1736 664
rect 1338 630 1355 653
tri 1355 630 1378 653 nw
tri 1696 630 1719 653 ne
rect 1719 630 1736 653
rect 1770 653 2168 664
rect 1770 630 1787 653
tri 1787 630 1810 653 nw
tri 2128 630 2151 653 ne
rect 2151 630 2168 653
rect 2202 630 2208 664
rect 756 621 1346 630
tri 1346 621 1355 630 nw
tri 1719 621 1728 630 ne
rect 1728 621 1776 630
rect 756 605 1344 621
tri 1344 619 1346 621 nw
rect 756 571 762 605
rect 796 571 1194 605
rect 1228 587 1344 605
rect 1228 571 1304 587
rect 756 559 1304 571
tri 1264 553 1270 559 ne
rect 1270 553 1304 559
rect 1338 553 1344 587
tri 1270 533 1290 553 ne
rect 1290 533 1344 553
tri 1290 525 1298 533 ne
tri 476 510 481 515 sw
rect 1298 510 1344 533
rect 214 481 481 510
tri 481 481 510 510 sw
rect 214 475 1270 481
rect 214 441 226 475
rect 260 441 303 475
rect 337 441 379 475
rect 413 441 455 475
rect 489 441 531 475
rect 565 441 607 475
rect 641 441 683 475
rect 717 441 759 475
rect 793 441 835 475
rect 869 441 911 475
rect 945 441 987 475
rect 1021 441 1063 475
rect 1097 441 1139 475
rect 1173 441 1270 475
rect 214 435 1270 441
tri 1128 433 1130 435 ne
rect 1130 433 1270 435
tri 1130 401 1162 433 ne
rect 269 155 351 164
rect 269 121 281 155
rect 315 121 351 155
rect 269 112 351 121
rect 403 112 415 164
rect 467 162 482 164
tri 482 162 484 164 sw
rect 467 161 484 162
tri 484 161 485 162 sw
rect 467 156 485 161
tri 485 156 490 161 sw
rect 467 122 490 156
tri 490 122 524 156 sw
rect 467 121 524 122
tri 524 121 525 122 sw
rect 467 118 525 121
tri 525 118 528 121 sw
rect 467 116 528 118
tri 528 116 530 118 sw
rect 467 115 530 116
tri 530 115 531 116 sw
rect 467 112 531 115
tri 531 112 534 115 sw
rect 603 113 609 165
rect 661 113 673 165
rect 725 113 762 165
rect 810 119 816 171
rect 868 119 880 171
rect 932 119 940 171
rect 810 115 940 119
rect 1001 119 1009 171
rect 1061 119 1073 171
rect 1125 119 1131 171
rect 1001 115 1131 119
tri 676 112 677 113 ne
rect 677 112 762 113
tri 468 89 491 112 ne
rect 491 89 534 112
tri 534 89 557 112 sw
tri 677 107 682 112 ne
rect 682 107 762 112
tri 682 89 700 107 ne
rect 700 89 762 107
tri 762 89 780 107 sw
tri 491 77 503 89 ne
rect 503 77 557 89
tri 557 77 569 89 sw
tri 700 79 710 89 ne
rect 710 77 780 89
tri 780 77 792 89 sw
rect 204 25 210 77
rect 262 25 274 77
rect 326 65 462 77
tri 503 74 506 77 ne
rect 506 74 569 77
tri 569 74 572 77 sw
rect 710 74 792 77
tri 792 74 795 77 sw
rect 326 31 422 65
rect 456 31 462 65
tri 506 61 519 74 ne
rect 519 73 572 74
tri 572 73 573 74 sw
rect 710 73 795 74
tri 795 73 796 74 sw
rect 519 61 573 73
tri 573 61 585 73 sw
rect 710 61 1102 73
tri 519 52 528 61 ne
rect 528 52 585 61
tri 585 52 594 61 sw
tri 528 40 540 52 ne
rect 540 40 678 52
rect 326 25 462 31
tri 540 28 552 40 ne
rect 552 28 678 40
rect 204 -6 253 25
tri 253 -6 284 25 nw
tri 382 -6 413 25 ne
rect 413 -6 462 25
tri 552 11 569 28 ne
rect 569 11 638 28
tri 598 -6 615 11 ne
rect 615 -6 638 11
rect 672 -6 678 28
rect 710 27 850 61
rect 884 27 1062 61
rect 1096 27 1102 61
rect 710 21 1102 27
tri 810 11 820 21 ne
rect 820 11 914 21
tri 914 11 924 21 nw
tri 1022 11 1032 21 ne
rect 1032 11 1102 21
tri 820 -3 834 11 ne
rect 834 -3 900 11
tri 900 -3 914 11 nw
tri 1032 -3 1046 11 ne
rect 1046 -3 1102 11
rect 204 -7 252 -6
tri 252 -7 253 -6 nw
tri 413 -7 414 -6 ne
rect 414 -7 462 -6
rect 204 -41 210 -7
rect 244 -41 250 -7
tri 250 -9 252 -7 nw
tri 414 -9 416 -7 ne
rect 204 -53 250 -41
rect 310 -44 356 -32
rect 310 -78 316 -44
rect 350 -78 356 -44
rect 416 -41 422 -7
rect 456 -41 462 -7
tri 615 -11 620 -6 ne
rect 620 -11 678 -6
tri 834 -11 842 -3 ne
rect 842 -11 892 -3
tri 892 -11 900 -3 nw
tri 1046 -11 1054 -3 ne
rect 1054 -11 1102 -3
tri 620 -23 632 -11 ne
rect 416 -53 462 -41
rect 522 -44 568 -32
rect 310 -116 356 -78
tri 286 -150 310 -126 se
rect 310 -150 316 -116
rect 350 -150 356 -116
rect 522 -78 528 -44
rect 562 -78 568 -44
rect 522 -116 568 -78
rect 632 -44 678 -11
tri 842 -13 844 -11 ne
rect 632 -78 638 -44
rect 672 -78 678 -44
rect 632 -90 678 -78
rect 738 -44 784 -32
rect 738 -78 744 -44
rect 778 -78 784 -44
rect 844 -45 850 -11
rect 884 -45 890 -11
tri 890 -13 892 -11 nw
tri 1054 -13 1056 -11 ne
rect 844 -57 890 -45
rect 950 -44 996 -32
tri 356 -150 380 -126 sw
tri 498 -150 522 -126 se
rect 522 -150 528 -116
rect 562 -150 568 -116
rect 738 -116 784 -78
tri 568 -150 592 -126 sw
tri 714 -150 738 -126 se
rect 738 -150 744 -116
rect 778 -150 784 -116
rect 950 -78 956 -44
rect 990 -78 996 -44
rect 1056 -45 1062 -11
rect 1096 -45 1102 -11
rect 1056 -57 1102 -45
rect 1162 -44 1270 433
rect 1298 476 1304 510
rect 1338 476 1344 510
rect 1298 433 1344 476
rect 1298 399 1304 433
rect 1338 399 1344 433
rect 1298 356 1344 399
rect 1298 322 1304 356
rect 1338 322 1344 356
rect 1298 279 1344 322
rect 1298 245 1304 279
rect 1338 245 1344 279
rect 1298 201 1344 245
rect 1298 167 1304 201
rect 1338 167 1344 201
rect 1298 123 1344 167
rect 1298 89 1304 123
rect 1338 89 1344 123
rect 1298 45 1344 89
rect 1298 11 1304 45
rect 1338 11 1344 45
rect 1298 -1 1344 11
rect 1511 615 1563 621
tri 1728 619 1730 621 ne
rect 1511 543 1563 563
rect 1511 471 1563 491
rect 1511 398 1563 419
rect 1511 325 1563 346
rect 1511 271 1520 273
rect 1554 271 1563 273
rect 1511 252 1563 271
rect 1511 194 1520 200
rect 1554 194 1563 200
rect 1511 151 1563 194
rect 1511 117 1520 151
rect 1554 117 1563 151
rect 1511 74 1563 117
rect 1511 40 1520 74
rect 1554 40 1563 74
rect 950 -116 996 -78
tri 784 -150 808 -126 sw
tri 926 -150 950 -126 se
rect 950 -150 956 -116
rect 990 -150 996 -116
rect 1162 -78 1168 -44
rect 1202 -78 1270 -44
rect 1162 -116 1270 -78
tri 996 -150 1020 -126 sw
tri 1138 -150 1162 -126 se
rect 1162 -150 1168 -116
rect 1202 -131 1270 -116
rect 1511 -3 1563 40
rect 1730 587 1776 621
tri 1776 619 1787 630 nw
tri 2151 619 2162 630 ne
rect 1730 553 1736 587
rect 1770 553 1776 587
rect 1730 510 1776 553
rect 2162 587 2208 630
rect 2162 553 2168 587
rect 2202 553 2208 587
rect 1730 476 1736 510
rect 1770 476 1776 510
rect 1730 433 1776 476
rect 1730 399 1736 433
rect 1770 399 1776 433
rect 1730 356 1776 399
rect 1730 322 1736 356
rect 1770 322 1776 356
rect 1730 279 1776 322
rect 1730 245 1736 279
rect 1770 245 1776 279
rect 1730 201 1776 245
rect 1730 167 1736 201
rect 1770 167 1776 201
rect 1730 123 1776 167
rect 1730 89 1736 123
rect 1770 89 1776 123
rect 1730 45 1776 89
rect 1730 11 1736 45
rect 1770 11 1776 45
rect 1730 -1 1776 11
rect 1946 521 1992 533
rect 1946 487 1952 521
rect 1986 487 1992 521
rect 1946 444 1992 487
rect 1946 410 1952 444
rect 1986 410 1992 444
rect 1946 367 1992 410
rect 1946 333 1952 367
rect 1986 333 1992 367
rect 1946 290 1992 333
rect 1946 256 1952 290
rect 1986 256 1992 290
rect 1946 213 1992 256
rect 1946 179 1952 213
rect 1986 179 1992 213
rect 1946 136 1992 179
rect 1946 102 1952 136
rect 1986 102 1992 136
rect 1946 59 1992 102
rect 1946 25 1952 59
rect 1986 25 1992 59
rect 1511 -37 1520 -3
rect 1554 -37 1563 -3
rect 1511 -80 1563 -37
rect 1511 -114 1520 -80
rect 1554 -114 1563 -80
rect 1511 -126 1563 -114
rect 1946 -19 1992 25
rect 2162 510 2208 553
rect 2162 476 2168 510
rect 2202 476 2208 510
rect 2162 433 2208 476
rect 2162 399 2168 433
rect 2202 399 2208 433
rect 2162 356 2208 399
rect 2162 322 2168 356
rect 2202 322 2208 356
rect 2162 279 2208 322
rect 2162 245 2168 279
rect 2202 245 2208 279
rect 2162 201 2208 245
rect 2162 167 2168 201
rect 2202 167 2208 201
rect 2162 123 2208 167
rect 2162 89 2168 123
rect 2202 89 2208 123
rect 2162 45 2208 89
rect 2162 11 2168 45
rect 2202 11 2208 45
rect 2162 -1 2208 11
rect 2272 741 2318 753
rect 2272 707 2278 741
rect 2312 707 2318 741
rect 2272 665 2318 707
rect 2272 631 2278 665
rect 2312 631 2318 665
rect 2272 589 2318 631
rect 2272 555 2278 589
rect 2312 555 2318 589
rect 2272 513 2318 555
rect 2272 479 2278 513
rect 2312 479 2318 513
rect 2272 437 2318 479
rect 2272 403 2278 437
rect 2312 403 2318 437
rect 2272 361 2318 403
rect 2272 327 2278 361
rect 2312 327 2318 361
rect 2272 285 2318 327
rect 2272 251 2278 285
rect 2312 251 2318 285
rect 2272 209 2318 251
rect 2272 175 2278 209
rect 2312 175 2318 209
rect 2272 133 2318 175
rect 2272 99 2278 133
rect 2312 99 2318 133
rect 2272 56 2318 99
rect 2272 22 2278 56
rect 2312 22 2318 56
rect 1946 -53 1952 -19
rect 1986 -53 1992 -19
rect 1946 -97 1992 -53
tri 1270 -131 1275 -126 sw
tri 1941 -131 1946 -126 se
rect 1946 -131 1952 -97
rect 1986 -131 1992 -97
rect 2272 -21 2318 22
rect 2272 -55 2278 -21
rect 2312 -55 2318 -21
rect 2272 -98 2318 -55
rect 1202 -132 1275 -131
tri 1275 -132 1276 -131 sw
tri 1940 -132 1941 -131 se
rect 1941 -132 1992 -131
tri 1992 -132 1998 -126 sw
tri 2266 -132 2272 -126 se
rect 2272 -132 2278 -98
rect 2312 -132 2318 -98
rect 2488 741 2534 834
rect 2488 707 2494 741
rect 2528 707 2534 741
rect 2488 665 2534 707
rect 2488 631 2494 665
rect 2528 631 2534 665
rect 2488 589 2534 631
rect 2488 555 2494 589
rect 2528 555 2534 589
rect 2488 513 2534 555
rect 2488 479 2494 513
rect 2528 479 2534 513
rect 2488 437 2534 479
rect 2488 403 2494 437
rect 2528 403 2534 437
rect 2488 361 2534 403
rect 2488 327 2494 361
rect 2528 327 2534 361
rect 2488 285 2534 327
rect 2488 251 2494 285
rect 2528 251 2534 285
rect 2488 209 2534 251
rect 2488 175 2494 209
rect 2528 175 2534 209
rect 2488 133 2534 175
rect 2488 99 2494 133
rect 2528 99 2534 133
rect 2488 56 2534 99
rect 2488 22 2494 56
rect 2528 22 2534 56
rect 2488 -21 2534 22
rect 2488 -55 2494 -21
rect 2528 -55 2534 -21
rect 2488 -98 2534 -55
tri 2318 -132 2324 -126 sw
tri 2482 -132 2488 -126 se
rect 2488 -132 2494 -98
rect 2528 -132 2534 -98
rect 1202 -150 1276 -132
tri 276 -160 286 -150 se
rect 286 -160 380 -150
tri 380 -160 390 -150 sw
tri 488 -160 498 -150 se
rect 498 -160 592 -150
tri 592 -160 602 -150 sw
tri 704 -160 714 -150 se
rect 714 -160 808 -150
tri 808 -160 818 -150 sw
tri 916 -160 926 -150 se
rect 926 -160 1020 -150
tri 1020 -160 1030 -150 sw
tri 1128 -160 1138 -150 se
rect 1138 -160 1276 -150
tri 1276 -160 1304 -132 sw
tri 1912 -160 1940 -132 se
rect 1940 -160 1998 -132
tri 1998 -160 2026 -132 sw
tri 2238 -160 2266 -132 se
rect 2266 -160 2324 -132
tri 2324 -160 2352 -132 sw
tri 2454 -160 2482 -132 se
rect 2482 -160 2534 -132
tri 2534 -160 2568 -126 sw
rect 114 -175 2586 -160
rect 114 -209 1952 -175
rect 1986 -209 2278 -175
rect 2312 -209 2494 -175
rect 2528 -209 2586 -175
rect 114 -281 2586 -209
rect 114 -315 172 -281
rect 206 -315 246 -281
rect 280 -315 320 -281
rect 354 -315 394 -281
rect 428 -315 468 -281
rect 502 -315 542 -281
rect 576 -315 616 -281
rect 650 -315 690 -281
rect 724 -315 764 -281
rect 798 -315 838 -281
rect 872 -315 912 -281
rect 946 -315 986 -281
rect 1020 -315 1060 -281
rect 1094 -315 1134 -281
rect 1168 -315 1208 -281
rect 1242 -315 1282 -281
rect 1316 -315 1355 -281
rect 1389 -315 1428 -281
rect 1462 -315 1501 -281
rect 1535 -315 1574 -281
rect 1608 -315 1647 -281
rect 1681 -315 1720 -281
rect 1754 -315 1793 -281
rect 1827 -315 1866 -281
rect 1900 -315 1939 -281
rect 1973 -315 2012 -281
rect 2046 -315 2085 -281
rect 2119 -315 2158 -281
rect 2192 -315 2231 -281
rect 2265 -315 2304 -281
rect 2338 -315 2377 -281
rect 2411 -315 2450 -281
rect 2484 -315 2586 -281
rect 114 -575 2586 -315
<< via1 >>
rect 671 3544 673 3577
rect 673 3544 707 3577
rect 707 3544 723 3577
rect 768 3544 784 3577
rect 784 3544 820 3577
rect 865 3544 904 3577
rect 904 3544 917 3577
rect 962 3544 981 3577
rect 981 3544 1014 3577
rect 1059 3544 1092 3577
rect 1092 3544 1111 3577
rect 1156 3544 1169 3577
rect 1169 3544 1208 3577
rect 671 3525 723 3544
rect 768 3525 820 3544
rect 865 3525 917 3544
rect 962 3525 1014 3544
rect 1059 3525 1111 3544
rect 1156 3525 1208 3544
rect 448 3425 500 3434
rect 448 3391 452 3425
rect 452 3391 486 3425
rect 486 3391 500 3425
rect 448 3382 500 3391
rect 512 3425 564 3434
rect 512 3391 524 3425
rect 524 3391 558 3425
rect 558 3391 564 3425
rect 512 3382 564 3391
rect 1248 3408 1300 3460
rect 1312 3454 1364 3460
rect 1312 3420 1330 3454
rect 1330 3420 1364 3454
rect 1312 3408 1364 3420
rect 1410 3480 1462 3488
rect 1410 3446 1414 3480
rect 1414 3446 1448 3480
rect 1448 3446 1462 3480
rect 1410 3436 1462 3446
rect 1474 3480 1526 3488
rect 1474 3446 1486 3480
rect 1486 3446 1520 3480
rect 1520 3446 1526 3480
rect 1474 3436 1526 3446
rect 1683 3534 1799 3639
rect 1683 3523 1694 3534
rect 1694 3523 1728 3534
rect 1728 3523 1799 3534
rect 1707 3390 1759 3412
rect 1707 3360 1728 3390
rect 1728 3360 1759 3390
rect 1707 3318 1759 3329
rect 1707 3284 1728 3318
rect 1728 3284 1759 3318
rect 1707 3277 1759 3284
rect 1032 3264 1084 3273
rect 1096 3264 1148 3273
rect 1032 3230 1061 3264
rect 1061 3230 1084 3264
rect 1096 3230 1140 3264
rect 1140 3230 1148 3264
rect 1032 3221 1084 3230
rect 1096 3221 1148 3230
rect 1707 3212 1728 3246
rect 1728 3212 1759 3246
rect 1707 3194 1759 3212
rect 444 3105 496 3114
rect 444 3071 450 3105
rect 450 3071 484 3105
rect 484 3071 496 3105
rect 444 3062 496 3071
rect 508 3105 560 3114
rect 508 3071 522 3105
rect 522 3071 556 3105
rect 556 3071 560 3105
rect 508 3062 560 3071
rect 1707 3140 1728 3163
rect 1728 3140 1759 3163
rect 1707 3111 1759 3140
rect 1707 3068 1728 3080
rect 1728 3068 1759 3080
rect 876 3052 928 3061
rect 940 3052 992 3061
rect 876 3018 903 3052
rect 903 3018 928 3052
rect 940 3018 982 3052
rect 982 3018 992 3052
rect 876 3009 928 3018
rect 940 3009 992 3018
rect 1707 3029 1759 3068
rect 1707 3028 1728 3029
rect 1728 3028 1759 3029
rect 1707 2995 1728 2997
rect 1728 2995 1759 2997
rect 1707 2956 1759 2995
rect 708 2942 760 2951
rect 772 2942 824 2951
rect 708 2908 745 2942
rect 745 2908 760 2942
rect 772 2908 779 2942
rect 779 2908 824 2942
rect 708 2899 760 2908
rect 772 2899 824 2908
rect 1707 2945 1728 2956
rect 1728 2945 1759 2956
rect 448 2891 500 2899
rect 448 2857 452 2891
rect 452 2857 486 2891
rect 486 2857 500 2891
rect 448 2847 500 2857
rect 512 2891 564 2899
rect 512 2857 524 2891
rect 524 2857 558 2891
rect 558 2857 564 2891
rect 512 2847 564 2857
rect 1707 2883 1759 2914
rect 1707 2862 1728 2883
rect 1728 2862 1759 2883
rect 1707 2810 1759 2831
rect 1707 2779 1728 2810
rect 1728 2779 1759 2810
rect 521 2649 530 2677
rect 530 2649 564 2677
rect 564 2649 573 2677
rect 521 2625 573 2649
rect 521 2601 573 2613
rect 521 2567 530 2601
rect 530 2567 564 2601
rect 564 2567 573 2601
rect 521 2561 573 2567
rect 1180 2730 1232 2739
rect 1244 2730 1296 2739
rect 1180 2696 1219 2730
rect 1219 2696 1232 2730
rect 1244 2696 1253 2730
rect 1253 2696 1296 2730
rect 1180 2687 1232 2696
rect 1244 2687 1296 2696
rect 1707 2737 1759 2748
rect 1707 2703 1728 2737
rect 1728 2703 1759 2737
rect 1707 2696 1759 2703
rect 1707 2664 1759 2665
rect 1707 2630 1728 2664
rect 1728 2630 1759 2664
rect 1707 2613 1759 2630
rect 1707 2530 1759 2582
rect 1180 2518 1232 2527
rect 1244 2518 1296 2527
rect 1180 2484 1219 2518
rect 1219 2484 1232 2518
rect 1244 2484 1253 2518
rect 1253 2484 1296 2518
rect 1180 2475 1232 2484
rect 1244 2475 1296 2484
rect 1707 2446 1759 2498
rect 527 2266 579 2318
rect 591 2266 643 2318
rect 788 2266 840 2318
rect 852 2266 904 2318
rect 480 2182 532 2234
rect 544 2182 596 2234
rect 1822 2182 1874 2234
rect 1886 2182 1938 2234
rect 1180 2002 1232 2011
rect 1244 2002 1296 2011
rect 1180 1968 1195 2002
rect 1195 1968 1232 2002
rect 1244 1968 1272 2002
rect 1272 1968 1296 2002
rect 1180 1959 1232 1968
rect 1244 1959 1296 1968
rect 1707 1997 1759 2003
rect 1707 1963 1716 1997
rect 1716 1963 1750 1997
rect 1750 1963 1759 1997
rect 1707 1951 1759 1963
rect 550 1915 602 1921
rect 550 1881 560 1915
rect 560 1881 594 1915
rect 594 1881 602 1915
rect 550 1869 602 1881
rect 1707 1925 1759 1937
rect 1707 1891 1716 1925
rect 1716 1891 1750 1925
rect 1750 1891 1759 1925
rect 1707 1885 1759 1891
rect 550 1823 602 1857
rect 550 1805 560 1823
rect 560 1805 594 1823
rect 594 1805 602 1823
rect 866 1791 918 1843
rect 1330 1816 1382 1868
rect 1707 1853 1759 1871
rect 1707 1819 1716 1853
rect 1716 1819 1750 1853
rect 1750 1819 1759 1853
rect 1330 1786 1382 1804
rect 1496 1786 1548 1794
rect 1560 1786 1612 1794
rect 866 1752 889 1779
rect 889 1752 918 1779
rect 1330 1752 1356 1786
rect 1356 1752 1382 1786
rect 1496 1752 1510 1786
rect 1510 1752 1548 1786
rect 1560 1752 1587 1786
rect 1587 1752 1612 1786
rect 866 1727 918 1752
rect 1496 1742 1548 1752
rect 1560 1742 1612 1752
rect 1707 1781 1759 1805
rect 1707 1753 1716 1781
rect 1716 1753 1750 1781
rect 1750 1753 1759 1781
rect 1707 1709 1759 1739
rect 1707 1687 1716 1709
rect 1716 1687 1750 1709
rect 1750 1687 1759 1709
rect 1707 1636 1759 1672
rect 1707 1620 1716 1636
rect 1716 1620 1750 1636
rect 1750 1620 1759 1636
rect 1707 1602 1716 1605
rect 1716 1602 1750 1605
rect 1750 1602 1759 1605
rect 1180 1570 1232 1579
rect 1180 1536 1201 1570
rect 1201 1536 1232 1570
rect 1180 1527 1232 1536
rect 1244 1570 1296 1579
rect 1244 1536 1245 1570
rect 1245 1536 1279 1570
rect 1279 1536 1296 1570
rect 1244 1527 1296 1536
rect 1707 1563 1759 1602
rect 1707 1553 1716 1563
rect 1716 1553 1750 1563
rect 1750 1553 1759 1563
rect 341 1468 393 1520
rect 341 1404 393 1456
rect 533 1398 585 1450
rect 597 1398 649 1450
rect 1340 1398 1392 1450
rect 1404 1398 1456 1450
rect 427 1318 479 1370
rect 491 1318 543 1370
rect 952 1318 1004 1370
rect 1016 1318 1068 1370
rect 210 1238 262 1290
rect 274 1238 326 1290
rect 1108 1238 1160 1290
rect 1172 1238 1224 1290
rect 788 1090 840 1142
rect 852 1090 904 1142
rect 1109 1090 1161 1142
rect 1173 1090 1225 1142
rect 872 877 924 886
rect 872 843 905 877
rect 905 843 924 877
rect 872 834 924 843
rect 936 877 988 886
rect 936 843 950 877
rect 950 843 984 877
rect 984 843 988 877
rect 936 834 988 843
rect 1822 877 1874 886
rect 1822 843 1850 877
rect 1850 843 1874 877
rect 1822 834 1874 843
rect 1886 877 1938 886
rect 1886 843 1890 877
rect 1890 843 1924 877
rect 1924 843 1938 877
rect 1886 834 1938 843
rect 708 732 760 784
rect 772 732 824 784
rect 351 155 403 164
rect 351 121 353 155
rect 353 121 387 155
rect 387 121 403 155
rect 351 112 403 121
rect 415 112 467 164
rect 609 156 661 165
rect 609 122 615 156
rect 615 122 649 156
rect 649 122 661 156
rect 609 113 661 122
rect 673 156 725 165
rect 673 122 687 156
rect 687 122 721 156
rect 721 122 725 156
rect 673 113 725 122
rect 816 155 868 171
rect 816 121 822 155
rect 822 121 856 155
rect 856 121 868 155
rect 816 119 868 121
rect 880 155 932 171
rect 880 121 894 155
rect 894 121 928 155
rect 928 121 932 155
rect 880 119 932 121
rect 1009 155 1061 171
rect 1009 121 1013 155
rect 1013 121 1047 155
rect 1047 121 1061 155
rect 1009 119 1061 121
rect 1073 155 1125 171
rect 1073 121 1085 155
rect 1085 121 1119 155
rect 1119 121 1125 155
rect 1073 119 1125 121
rect 210 65 262 77
rect 210 31 244 65
rect 244 31 262 65
rect 210 25 262 31
rect 274 25 326 77
rect 1511 609 1563 615
rect 1511 575 1520 609
rect 1520 575 1554 609
rect 1554 575 1563 609
rect 1511 563 1563 575
rect 1511 533 1563 543
rect 1511 499 1520 533
rect 1520 499 1554 533
rect 1554 499 1563 533
rect 1511 491 1563 499
rect 1511 457 1563 471
rect 1511 423 1520 457
rect 1520 423 1554 457
rect 1554 423 1563 457
rect 1511 419 1563 423
rect 1511 381 1563 398
rect 1511 347 1520 381
rect 1520 347 1554 381
rect 1554 347 1563 381
rect 1511 346 1563 347
rect 1511 305 1563 325
rect 1511 273 1520 305
rect 1520 273 1554 305
rect 1554 273 1563 305
rect 1511 228 1563 252
rect 1511 200 1520 228
rect 1520 200 1554 228
rect 1554 200 1563 228
<< metal2 >>
rect 665 3639 1799 3645
rect 665 3577 1683 3639
rect 665 3525 671 3577
rect 723 3525 768 3577
rect 820 3525 865 3577
rect 917 3525 962 3577
rect 1014 3525 1059 3577
rect 1111 3525 1156 3577
rect 1208 3525 1683 3577
rect 665 3523 1683 3525
rect 665 3517 1799 3523
rect 437 3382 448 3434
rect 500 3382 512 3434
rect 564 3382 658 3434
rect 1242 3408 1248 3460
rect 1300 3408 1312 3460
rect 1364 3408 1370 3460
rect 1404 3436 1410 3488
rect 1462 3436 1474 3488
rect 1526 3436 1532 3488
tri 1446 3434 1448 3436 ne
rect 1448 3434 1532 3436
tri 1448 3412 1470 3434 ne
rect 1470 3412 1532 3434
tri 1470 3408 1474 3412 ne
rect 1474 3408 1532 3412
tri 578 3360 600 3382 ne
rect 600 3360 658 3382
tri 1252 3376 1284 3408 ne
rect 1284 3376 1338 3408
tri 1338 3376 1370 3408 nw
tri 1474 3402 1480 3408 ne
tri 1284 3374 1286 3376 ne
tri 600 3348 612 3360 ne
tri 348 3062 400 3114 se
rect 400 3062 444 3114
rect 496 3062 508 3114
rect 560 3062 566 3114
tri 606 3062 612 3068 se
rect 612 3062 658 3360
rect 1026 3221 1032 3273
rect 1084 3221 1096 3273
rect 1148 3221 1154 3273
rect 1286 3221 1338 3376
tri 1338 3221 1353 3236 sw
tri 1026 3199 1048 3221 ne
tri 347 3061 348 3062 se
rect 348 3061 421 3062
tri 421 3061 422 3062 nw
tri 605 3061 606 3062 se
rect 606 3061 658 3062
rect 1048 3194 1107 3221
tri 1107 3194 1134 3221 nw
rect 1286 3214 1353 3221
tri 1286 3194 1306 3214 ne
rect 1306 3194 1353 3214
tri 1353 3194 1380 3221 sw
tri 341 3055 347 3061 se
rect 347 3055 415 3061
tri 415 3055 421 3061 nw
tri 599 3055 605 3061 se
rect 605 3055 658 3061
rect 341 1520 393 3055
tri 393 3033 415 3055 nw
tri 577 3033 599 3055 se
rect 599 3048 658 3055
rect 599 3033 619 3048
tri 553 3009 577 3033 se
rect 577 3009 619 3033
tri 619 3009 658 3048 nw
rect 870 3009 876 3061
rect 928 3009 940 3061
rect 992 3009 998 3061
tri 546 3002 553 3009 se
rect 553 3002 612 3009
tri 612 3002 619 3009 nw
tri 912 3002 919 3009 ne
rect 919 3002 998 3009
tri 541 2997 546 3002 se
rect 546 2997 607 3002
tri 607 2997 612 3002 nw
tri 919 2997 924 3002 ne
rect 924 2997 998 3002
tri 524 2980 541 2997 se
rect 541 2980 590 2997
tri 590 2980 607 2997 nw
tri 924 2980 941 2997 ne
rect 941 2980 998 2997
tri 490 2899 524 2933 se
rect 524 2899 570 2980
tri 570 2960 590 2980 nw
tri 941 2975 946 2980 ne
rect 442 2847 448 2899
rect 500 2847 512 2899
rect 564 2847 570 2899
rect 702 2899 708 2951
rect 760 2899 772 2951
rect 824 2899 830 2951
rect 521 2677 573 2683
rect 521 2613 573 2625
rect 521 2318 573 2561
tri 573 2318 607 2352 sw
rect 521 2266 527 2318
rect 579 2266 591 2318
rect 643 2266 649 2318
rect 474 2182 480 2234
rect 532 2182 544 2234
rect 596 2182 602 2234
tri 516 2148 550 2182 ne
rect 550 1921 602 2182
rect 550 1857 602 1869
rect 550 1799 602 1805
rect 341 1456 393 1468
rect 341 1398 393 1404
rect 527 1398 533 1450
rect 585 1398 597 1450
rect 649 1398 655 1450
tri 569 1370 597 1398 ne
rect 597 1370 655 1398
rect 421 1318 427 1370
rect 479 1318 491 1370
rect 543 1318 549 1370
tri 597 1364 603 1370 ne
rect 421 1290 479 1318
tri 479 1290 507 1318 nw
rect 204 1238 210 1290
rect 262 1238 274 1290
rect 326 1238 332 1290
rect 204 77 256 1238
tri 256 1204 290 1238 nw
tri 394 171 421 198 se
rect 421 171 473 1290
tri 473 1284 479 1290 nw
tri 388 165 394 171 se
rect 394 165 473 171
tri 387 164 388 165 se
rect 388 164 473 165
rect 345 112 351 164
rect 403 112 415 164
rect 467 112 473 164
rect 603 194 655 1370
rect 702 784 754 2899
tri 754 2865 788 2899 nw
rect 782 2266 788 2318
rect 840 2266 852 2318
rect 904 2266 910 2318
rect 782 2234 836 2266
tri 836 2234 868 2266 nw
rect 782 1142 834 2234
tri 834 2232 836 2234 nw
rect 866 1843 918 1849
rect 866 1779 918 1791
rect 866 1241 918 1727
rect 946 1398 998 2980
rect 1048 1478 1100 3194
tri 1100 3187 1107 3194 nw
tri 1306 3192 1308 3194 ne
rect 1308 3192 1380 3194
tri 1380 3192 1382 3194 sw
tri 1308 3187 1313 3192 ne
rect 1313 3187 1382 3192
tri 1313 3170 1330 3187 ne
rect 1174 2687 1180 2739
rect 1232 2687 1244 2739
rect 1296 2687 1302 2739
rect 1174 2527 1302 2687
rect 1174 2475 1180 2527
rect 1232 2475 1244 2527
rect 1296 2475 1302 2527
rect 1174 2011 1302 2475
rect 1174 1959 1180 2011
rect 1232 1959 1244 2011
rect 1296 1959 1302 2011
rect 1174 1579 1302 1959
rect 1330 1868 1382 3187
rect 1330 1804 1382 1816
rect 1330 1746 1382 1752
tri 1410 2112 1480 2182 se
rect 1480 2160 1532 3408
rect 1480 2112 1484 2160
tri 1484 2112 1532 2160 nw
rect 1707 3412 1759 3418
rect 1707 3329 1759 3360
rect 1707 3246 1759 3277
rect 1707 3163 1759 3194
rect 1707 3080 1759 3111
rect 1707 2997 1759 3028
rect 1707 2914 1759 2945
rect 1707 2831 1759 2862
rect 1707 2748 1759 2779
rect 1707 2665 1759 2696
rect 1707 2582 1759 2613
rect 1707 2498 1759 2530
rect 1174 1527 1180 1579
rect 1232 1527 1244 1579
rect 1296 1527 1302 1579
tri 1048 1450 1076 1478 ne
rect 1076 1450 1100 1478
tri 1100 1450 1150 1500 sw
tri 1376 1450 1410 1484 se
rect 1410 1450 1462 2112
tri 1462 2090 1484 2112 nw
rect 1707 2003 1759 2446
rect 1816 2182 1822 2234
rect 1874 2182 1886 2234
rect 1938 2182 1944 2234
tri 1858 2148 1892 2182 ne
rect 1707 1937 1759 1951
rect 1707 1871 1759 1885
rect 1707 1805 1759 1819
tri 1076 1446 1080 1450 ne
rect 1080 1446 1150 1450
tri 1150 1446 1154 1450 sw
tri 1080 1426 1100 1446 ne
rect 1100 1426 1154 1446
tri 1100 1424 1102 1426 ne
tri 998 1398 1004 1404 sw
rect 946 1370 1004 1398
tri 1004 1370 1032 1398 sw
rect 946 1318 952 1370
rect 1004 1318 1016 1370
rect 1068 1318 1074 1370
rect 1102 1318 1154 1426
rect 1334 1398 1340 1450
rect 1392 1398 1404 1450
rect 1456 1398 1462 1450
rect 1490 1742 1496 1794
rect 1548 1742 1560 1794
rect 1612 1742 1618 1794
tri 1154 1318 1160 1324 sw
rect 1102 1290 1160 1318
tri 1160 1290 1188 1318 sw
tri 918 1241 952 1275 sw
rect 866 1189 1050 1241
rect 1102 1238 1108 1290
rect 1160 1238 1172 1290
rect 1224 1238 1230 1290
tri 964 1181 972 1189 ne
rect 972 1181 1050 1189
tri 834 1142 873 1181 sw
tri 972 1155 998 1181 ne
rect 782 1090 788 1142
rect 840 1090 852 1142
rect 904 1090 910 1142
tri 964 886 998 920 se
rect 998 886 1050 1181
rect 866 834 872 886
rect 924 834 936 886
rect 988 834 1050 886
rect 1103 1090 1109 1142
rect 1161 1090 1173 1142
rect 1225 1090 1231 1142
rect 866 818 936 834
tri 936 818 952 834 nw
tri 754 784 788 818 sw
rect 702 732 708 784
rect 760 732 772 784
rect 824 732 830 784
tri 861 200 866 205 se
rect 866 200 918 818
tri 918 800 936 818 nw
tri 1098 200 1103 205 se
rect 1103 200 1155 1090
tri 1155 1061 1184 1090 nw
tri 860 199 861 200 se
rect 861 199 918 200
tri 655 194 660 199 sw
tri 855 194 860 199 se
rect 860 194 918 199
tri 1092 194 1098 200 se
rect 1098 194 1155 200
rect 1490 615 1618 1742
rect 1707 1739 1759 1753
rect 1707 1672 1759 1687
rect 1707 1605 1759 1620
rect 1707 1547 1759 1553
tri 1858 886 1892 920 se
rect 1892 886 1944 2182
rect 1816 834 1822 886
rect 1874 834 1886 886
rect 1938 834 1944 886
rect 1490 563 1511 615
rect 1563 563 1618 615
rect 1490 543 1618 563
rect 1490 491 1511 543
rect 1563 491 1618 543
rect 1490 471 1618 491
rect 1490 419 1511 471
rect 1563 419 1618 471
rect 1490 398 1618 419
rect 1490 346 1511 398
rect 1563 346 1618 398
rect 1490 325 1618 346
rect 1490 273 1511 325
rect 1563 273 1618 325
rect 1490 252 1618 273
rect 1490 200 1511 252
rect 1563 200 1618 252
rect 1490 194 1618 200
rect 603 171 660 194
tri 660 171 683 194 sw
tri 832 171 855 194 se
rect 855 171 918 194
tri 1089 191 1092 194 se
rect 1092 191 1155 194
tri 918 171 938 191 sw
tri 1069 171 1089 191 se
rect 1089 171 1155 191
rect 603 165 683 171
tri 683 165 689 171 sw
rect 603 113 609 165
rect 661 113 673 165
rect 725 113 731 165
rect 810 119 816 171
rect 868 119 880 171
rect 932 119 938 171
rect 1003 119 1009 171
rect 1061 119 1073 171
rect 1125 119 1155 171
tri 256 77 290 111 sw
rect 204 25 210 77
rect 262 25 274 77
rect 326 25 332 77
use sky130_fd_pr__nfet_01v8__example_5595914180825  sky130_fd_pr__nfet_01v8__example_5595914180825_0
timestamp 1683767628
transform 1 0 683 0 -1 73
box -1 0 51 1
use sky130_fd_pr__nfet_01v8__example_55959141808527  sky130_fd_pr__nfet_01v8__example_55959141808527_0
timestamp 1683767628
transform -1 0 1183 0 1 595
box -1 0 593 1
use sky130_fd_pr__nfet_01v8__example_55959141808535  sky130_fd_pr__nfet_01v8__example_55959141808535_0
timestamp 1683767628
transform 1 0 1349 0 1 -205
box -1 0 377 1
use sky130_fd_pr__nfet_01v8__example_55959141808535  sky130_fd_pr__nfet_01v8__example_55959141808535_1
timestamp 1683767628
transform 1 0 1781 0 1 -205
box -1 0 377 1
use sky130_fd_pr__nfet_01v8__example_55959141808601  sky130_fd_pr__nfet_01v8__example_55959141808601_0
timestamp 1683767628
transform 1 0 255 0 -1 73
box -1 0 263 1
use sky130_fd_pr__nfet_01v8__example_55959141808602  sky130_fd_pr__nfet_01v8__example_55959141808602_0
timestamp 1683767628
transform 1 0 789 0 -1 73
box -1 0 157 1
use sky130_fd_pr__nfet_01v8__example_55959141808602  sky130_fd_pr__nfet_01v8__example_55959141808602_1
timestamp 1683767628
transform 1 0 1001 0 -1 73
box -1 0 157 1
use sky130_fd_pr__nfet_01v8__example_55959141808603  sky130_fd_pr__nfet_01v8__example_55959141808603_0
timestamp 1683767628
transform -1 0 425 0 1 595
box -1 0 161 1
use sky130_fd_pr__nfet_01v8__example_55959141808604  sky130_fd_pr__nfet_01v8__example_55959141808604_0
timestamp 1683767628
transform 1 0 2323 0 1 -205
box -1 0 161 1
use sky130_fd_pr__pfet_01v8__example_55959141808540  sky130_fd_pr__pfet_01v8__example_55959141808540_0
timestamp 1683767628
transform 0 1 642 -1 0 1957
box -1 0 377 1
use sky130_fd_pr__pfet_01v8__example_55959141808596  sky130_fd_pr__pfet_01v8__example_55959141808596_0
timestamp 1683767628
transform 0 -1 1612 1 0 2847
box -1 0 51 1
use sky130_fd_pr__pfet_01v8__example_55959141808596  sky130_fd_pr__pfet_01v8__example_55959141808596_1
timestamp 1683767628
transform 0 -1 1612 -1 0 3113
box -1 0 51 1
use sky130_fd_pr__pfet_01v8__example_55959141808596  sky130_fd_pr__pfet_01v8__example_55959141808596_2
timestamp 1683767628
transform 0 -1 1612 -1 0 3219
box -1 0 51 1
use sky130_fd_pr__pfet_01v8__example_55959141808598  sky130_fd_pr__pfet_01v8__example_55959141808598_0
timestamp 1683767628
transform 0 -1 1212 1 0 3385
box -1 0 51 1
use sky130_fd_pr__pfet_01v8__example_55959141808605  sky130_fd_pr__pfet_01v8__example_55959141808605_0
timestamp 1683767628
transform 0 -1 1612 1 0 3385
box -1 0 157 1
use sky130_fd_pr__pfet_01v8__example_55959141808606  sky130_fd_pr__pfet_01v8__example_55959141808606_0
timestamp 1683767628
transform 0 -1 1612 -1 0 2791
box -1 0 263 1
<< labels >>
flabel metal1 s 625 2192 692 2229 3 FreeSans 200 0 0 0 IN_H
port 1 nsew
flabel metal1 s 481 2271 560 2309 3 FreeSans 200 0 0 0 MODE_VCCHIB_LV_N
port 2 nsew
flabel metal1 s 1622 2760 1781 3015 3 FreeSans 200 0 0 0 VCCHIB
port 3 nsew
flabel metal1 s 1194 -552 1780 -375 3 FreeSans 200 0 0 0 VSSD
port 4 nsew
flabel metal1 s 354 1251 412 1281 3 FreeSans 200 0 0 0 OUT
port 5 nsew
flabel metal1 s 561 1323 624 1360 3 FreeSans 200 0 0 0 OUT_N
port 6 nsew
<< properties >>
string GDS_END 3593004
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3527840
<< end >>
