magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 1 21 1165 203
rect 29 -17 63 21
<< scnmos >>
rect 82 47 112 177
rect 166 47 196 177
rect 250 47 280 177
rect 334 47 364 177
rect 522 47 552 177
rect 606 47 636 177
rect 690 47 720 177
rect 785 47 815 177
rect 973 47 1003 177
rect 1057 47 1087 177
<< scpmoshvt >>
rect 82 297 112 497
rect 166 297 196 497
rect 250 297 280 497
rect 334 297 364 497
rect 522 297 552 497
rect 606 297 636 497
rect 690 297 720 497
rect 785 297 815 497
rect 973 297 1003 497
rect 1057 297 1087 497
<< ndiff >>
rect 27 95 82 177
rect 27 61 38 95
rect 72 61 82 95
rect 27 47 82 61
rect 112 163 166 177
rect 112 129 122 163
rect 156 129 166 163
rect 112 95 166 129
rect 112 61 122 95
rect 156 61 166 95
rect 112 47 166 61
rect 196 95 250 177
rect 196 61 206 95
rect 240 61 250 95
rect 196 47 250 61
rect 280 163 334 177
rect 280 129 290 163
rect 324 129 334 163
rect 280 95 334 129
rect 280 61 290 95
rect 324 61 334 95
rect 280 47 334 61
rect 364 95 416 177
rect 364 61 374 95
rect 408 61 416 95
rect 364 47 416 61
rect 470 163 522 177
rect 470 129 478 163
rect 512 129 522 163
rect 470 95 522 129
rect 470 61 478 95
rect 512 61 522 95
rect 470 47 522 61
rect 552 95 606 177
rect 552 61 562 95
rect 596 61 606 95
rect 552 47 606 61
rect 636 125 690 177
rect 636 91 646 125
rect 680 91 690 125
rect 636 47 690 91
rect 720 163 785 177
rect 720 129 741 163
rect 775 129 785 163
rect 720 47 785 129
rect 815 95 867 177
rect 815 61 825 95
rect 859 61 867 95
rect 815 47 867 61
rect 921 95 973 177
rect 921 61 929 95
rect 963 61 973 95
rect 921 47 973 61
rect 1003 163 1057 177
rect 1003 129 1013 163
rect 1047 129 1057 163
rect 1003 47 1057 129
rect 1087 95 1139 177
rect 1087 61 1097 95
rect 1131 61 1139 95
rect 1087 47 1139 61
<< pdiff >>
rect 27 477 82 497
rect 27 443 38 477
rect 72 443 82 477
rect 27 297 82 443
rect 112 477 166 497
rect 112 443 122 477
rect 156 443 166 477
rect 112 297 166 443
rect 196 477 250 497
rect 196 443 206 477
rect 240 443 250 477
rect 196 297 250 443
rect 280 409 334 497
rect 280 375 290 409
rect 324 375 334 409
rect 280 297 334 375
rect 364 477 416 497
rect 364 443 374 477
rect 408 443 416 477
rect 364 297 416 443
rect 470 477 522 497
rect 470 443 478 477
rect 512 443 522 477
rect 470 409 522 443
rect 470 375 478 409
rect 512 375 522 409
rect 470 297 522 375
rect 552 477 606 497
rect 552 443 562 477
rect 596 443 606 477
rect 552 297 606 443
rect 636 477 690 497
rect 636 443 646 477
rect 680 443 690 477
rect 636 409 690 443
rect 636 375 646 409
rect 680 375 690 409
rect 636 297 690 375
rect 720 477 785 497
rect 720 443 741 477
rect 775 443 785 477
rect 720 297 785 443
rect 815 477 867 497
rect 815 443 825 477
rect 859 443 867 477
rect 815 409 867 443
rect 815 375 825 409
rect 859 375 867 409
rect 815 297 867 375
rect 921 477 973 497
rect 921 443 929 477
rect 963 443 973 477
rect 921 409 973 443
rect 921 375 929 409
rect 963 375 973 409
rect 921 297 973 375
rect 1003 409 1057 497
rect 1003 375 1013 409
rect 1047 375 1057 409
rect 1003 341 1057 375
rect 1003 307 1013 341
rect 1047 307 1057 341
rect 1003 297 1057 307
rect 1087 477 1143 497
rect 1087 443 1097 477
rect 1131 443 1143 477
rect 1087 409 1143 443
rect 1087 375 1097 409
rect 1131 375 1143 409
rect 1087 297 1143 375
<< ndiffc >>
rect 38 61 72 95
rect 122 129 156 163
rect 122 61 156 95
rect 206 61 240 95
rect 290 129 324 163
rect 290 61 324 95
rect 374 61 408 95
rect 478 129 512 163
rect 478 61 512 95
rect 562 61 596 95
rect 646 91 680 125
rect 741 129 775 163
rect 825 61 859 95
rect 929 61 963 95
rect 1013 129 1047 163
rect 1097 61 1131 95
<< pdiffc >>
rect 38 443 72 477
rect 122 443 156 477
rect 206 443 240 477
rect 290 375 324 409
rect 374 443 408 477
rect 478 443 512 477
rect 478 375 512 409
rect 562 443 596 477
rect 646 443 680 477
rect 646 375 680 409
rect 741 443 775 477
rect 825 443 859 477
rect 825 375 859 409
rect 929 443 963 477
rect 929 375 963 409
rect 1013 375 1047 409
rect 1013 307 1047 341
rect 1097 443 1131 477
rect 1097 375 1131 409
<< poly >>
rect 82 497 112 523
rect 166 497 196 523
rect 250 497 280 523
rect 334 497 364 523
rect 522 497 552 523
rect 606 497 636 523
rect 690 497 720 523
rect 785 497 815 523
rect 973 497 1003 523
rect 1057 497 1087 523
rect 82 265 112 297
rect 166 265 196 297
rect 250 265 280 297
rect 334 265 364 297
rect 522 265 552 297
rect 606 265 636 297
rect 690 265 720 297
rect 785 265 815 297
rect 82 249 196 265
rect 82 215 125 249
rect 159 215 196 249
rect 82 199 196 215
rect 248 249 364 265
rect 248 215 258 249
rect 292 215 364 249
rect 248 199 364 215
rect 518 249 640 265
rect 518 215 528 249
rect 562 215 596 249
rect 630 215 640 249
rect 518 199 640 215
rect 690 249 815 265
rect 690 215 700 249
rect 734 215 768 249
rect 802 215 815 249
rect 690 199 815 215
rect 82 177 112 199
rect 166 177 196 199
rect 250 177 280 199
rect 334 177 364 199
rect 522 177 552 199
rect 606 177 636 199
rect 690 177 720 199
rect 785 177 815 199
rect 973 265 1003 297
rect 1057 265 1087 297
rect 973 249 1087 265
rect 973 215 1005 249
rect 1039 215 1087 249
rect 973 199 1087 215
rect 973 177 1003 199
rect 1057 177 1087 199
rect 82 21 112 47
rect 166 21 196 47
rect 250 21 280 47
rect 334 21 364 47
rect 522 21 552 47
rect 606 21 636 47
rect 690 21 720 47
rect 785 21 815 47
rect 973 21 1003 47
rect 1057 21 1087 47
<< polycont >>
rect 125 215 159 249
rect 258 215 292 249
rect 528 215 562 249
rect 596 215 630 249
rect 700 215 734 249
rect 768 215 802 249
rect 1005 215 1039 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 24 477 80 493
rect 24 459 38 477
rect 24 427 29 459
rect 72 443 80 477
rect 63 427 80 443
rect 114 477 164 527
rect 114 443 122 477
rect 156 443 164 477
rect 114 427 164 443
rect 198 477 416 493
rect 198 443 206 477
rect 240 459 374 477
rect 198 427 213 443
rect 247 427 248 459
rect 366 443 374 459
rect 408 443 416 477
rect 366 427 416 443
rect 457 477 520 493
rect 457 443 478 477
rect 512 443 520 477
rect 457 425 520 443
rect 554 477 604 527
rect 554 443 562 477
rect 596 443 604 477
rect 554 427 604 443
rect 638 477 688 493
rect 638 443 646 477
rect 680 443 688 477
rect 282 409 332 425
rect 282 391 290 409
rect 24 375 290 391
rect 324 391 332 409
rect 478 409 520 425
rect 324 375 444 391
rect 24 357 444 375
rect 512 391 520 409
rect 638 409 688 443
rect 722 477 783 527
rect 722 443 741 477
rect 775 443 783 477
rect 722 427 783 443
rect 817 477 1139 493
rect 817 443 825 477
rect 859 443 929 477
rect 963 459 1097 477
rect 963 443 971 459
rect 638 391 646 409
rect 512 375 646 391
rect 680 391 688 409
rect 817 409 971 443
rect 1089 443 1097 459
rect 1131 443 1139 477
rect 817 391 825 409
rect 680 375 825 391
rect 859 375 929 409
rect 963 375 971 409
rect 478 357 971 375
rect 1005 409 1055 425
rect 1005 375 1013 409
rect 1047 375 1055 409
rect 24 181 58 357
rect 410 323 444 357
rect 1005 341 1055 375
rect 1089 409 1139 443
rect 1089 375 1097 409
rect 1131 375 1139 409
rect 1089 359 1139 375
rect 141 289 376 323
rect 410 289 957 323
rect 141 255 175 289
rect 342 255 376 289
rect 109 249 175 255
rect 109 215 125 249
rect 159 215 175 249
rect 209 221 213 255
rect 247 249 308 255
rect 247 221 258 249
rect 209 215 258 221
rect 292 215 308 249
rect 342 249 646 255
rect 342 215 528 249
rect 562 215 596 249
rect 630 215 646 249
rect 684 249 765 255
rect 799 249 818 255
rect 684 215 700 249
rect 734 221 765 249
rect 734 215 768 221
rect 802 215 818 249
rect 923 249 957 289
rect 1005 307 1013 341
rect 1047 325 1055 341
rect 1047 307 1179 325
rect 1005 283 1179 307
rect 923 215 1005 249
rect 1039 215 1055 249
rect 1097 181 1179 283
rect 24 163 340 181
rect 24 145 122 163
rect 106 129 122 145
rect 156 145 290 163
rect 156 129 172 145
rect 38 95 72 111
rect 38 17 72 61
rect 106 95 172 129
rect 274 129 290 145
rect 324 129 340 163
rect 106 61 122 95
rect 156 61 172 95
rect 106 51 172 61
rect 206 95 240 111
rect 206 17 240 61
rect 274 95 340 129
rect 462 163 680 181
rect 462 129 478 163
rect 512 145 680 163
rect 512 129 528 145
rect 274 61 290 95
rect 324 61 340 95
rect 274 51 340 61
rect 374 95 408 111
rect 374 17 408 61
rect 462 95 528 129
rect 630 125 680 145
rect 725 163 1179 181
rect 725 129 741 163
rect 775 145 1013 163
rect 775 129 791 145
rect 997 129 1013 145
rect 1047 145 1179 163
rect 1047 129 1063 145
rect 462 61 478 95
rect 512 61 528 95
rect 462 51 528 61
rect 562 95 596 111
rect 562 17 596 61
rect 630 91 646 125
rect 929 95 963 111
rect 680 91 825 95
rect 630 61 825 91
rect 859 61 876 95
rect 630 51 876 61
rect 929 17 963 61
rect 1097 95 1131 111
rect 1097 17 1131 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 443 38 459
rect 38 443 63 459
rect 29 425 63 443
rect 213 443 240 459
rect 240 443 247 459
rect 213 425 247 443
rect 213 221 247 255
rect 765 249 799 255
rect 765 221 768 249
rect 768 221 799 249
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 17 459 75 465
rect 17 425 29 459
rect 63 456 75 459
rect 201 459 259 465
rect 201 456 213 459
rect 63 428 213 456
rect 63 425 75 428
rect 17 419 75 425
rect 201 425 213 428
rect 247 425 259 459
rect 201 419 259 425
rect 201 255 259 261
rect 201 221 213 255
rect 247 252 259 255
rect 753 255 811 261
rect 753 252 765 255
rect 247 224 765 252
rect 247 221 259 224
rect 201 215 259 221
rect 753 221 765 224
rect 799 221 811 255
rect 753 215 811 221
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel locali s 1133 289 1167 323 0 FreeSans 400 0 0 0 X
port 7 nsew signal output
flabel locali s 765 221 799 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 213 289 247 323 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 xor2_2
rlabel locali s 684 215 818 255 1 B
port 2 nsew signal input
rlabel metal1 s 753 252 811 261 1 B
port 2 nsew signal input
rlabel metal1 s 753 215 811 224 1 B
port 2 nsew signal input
rlabel metal1 s 201 252 259 261 1 B
port 2 nsew signal input
rlabel metal1 s 201 224 811 252 1 B
port 2 nsew signal input
rlabel metal1 s 201 215 259 224 1 B
port 2 nsew signal input
rlabel metal1 s 0 -48 1196 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1196 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_END 646902
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 637824
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 2.720 5.980 2.720 
<< end >>
