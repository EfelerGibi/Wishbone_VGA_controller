magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< locali >>
rect 61039 65470 61073 65486
rect 61039 65420 61073 65436
<< viali >>
rect 61039 65436 61073 65470
<< metal1 >>
rect 61024 67361 61030 67413
rect 61082 67401 61088 67413
rect 64019 67401 64025 67413
rect 61082 67373 64025 67401
rect 61082 67361 61088 67373
rect 64019 67361 64025 67373
rect 64077 67361 64083 67413
rect 61024 65427 61030 65479
rect 61082 65427 61088 65479
<< via1 >>
rect 61030 67361 61082 67413
rect 64025 67361 64077 67413
rect 61030 65470 61082 65479
rect 61030 65436 61039 65470
rect 61039 65436 61073 65470
rect 61073 65436 61082 65470
rect 61030 65427 61082 65436
<< metal2 >>
rect 64037 67419 64065 68762
rect 61030 67413 61082 67419
rect 61030 67355 61082 67361
rect 64025 67413 64077 67419
rect 64025 67355 64077 67361
rect 61042 65485 61070 67355
rect 61030 65479 61082 65485
rect 61030 65421 61082 65427
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_0
timestamp 1683767628
transform 1 0 61027 0 1 65420
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_0
timestamp 1683767628
transform 1 0 64019 0 1 67355
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_1
timestamp 1683767628
transform 1 0 61024 0 1 65421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_2
timestamp 1683767628
transform 1 0 61024 0 1 67355
box 0 0 1 1
<< properties >>
string FIXED_BBOX 61024 65420 64083 68762
string GDS_END 7291198
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 7290450
<< end >>
