magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 1 201 1341 203
rect 1 23 1652 201
rect 1 21 197 23
rect 655 21 845 23
rect 1256 21 1652 23
rect 29 -17 63 21
<< locali >>
rect 17 288 73 493
rect 17 185 66 288
rect 17 70 69 185
rect 323 215 436 265
rect 1245 289 1361 323
rect 1245 199 1279 289
rect 1409 215 1491 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 107 443 174 527
rect 210 447 504 481
rect 645 447 711 527
rect 778 455 1397 489
rect 1479 455 1546 527
rect 210 409 244 447
rect 778 413 812 455
rect 107 375 244 409
rect 312 379 812 413
rect 107 265 141 375
rect 187 307 504 341
rect 100 199 141 265
rect 106 173 141 199
rect 106 139 221 173
rect 103 17 153 105
rect 187 85 221 139
rect 255 119 289 307
rect 470 265 504 307
rect 538 305 615 339
rect 559 275 615 305
rect 470 199 525 265
rect 349 159 425 181
rect 559 159 593 275
rect 649 241 683 379
rect 729 289 813 343
rect 349 125 593 159
rect 627 207 683 241
rect 627 91 661 207
rect 414 85 501 91
rect 187 51 501 85
rect 535 57 661 91
rect 695 17 729 173
rect 765 83 813 289
rect 849 119 883 421
rect 917 178 951 455
rect 1580 421 1639 493
rect 987 323 1070 409
rect 1177 387 1639 421
rect 987 289 1143 323
rect 990 199 1075 254
rect 917 165 959 178
rect 917 144 999 165
rect 925 131 999 144
rect 849 97 891 119
rect 849 53 931 97
rect 965 64 999 131
rect 1033 126 1075 199
rect 1109 85 1143 289
rect 1177 119 1211 387
rect 1542 375 1639 387
rect 1395 299 1559 341
rect 1525 265 1559 299
rect 1313 189 1375 255
rect 1525 199 1571 265
rect 1313 146 1354 189
rect 1525 181 1559 199
rect 1411 150 1559 181
rect 1403 147 1559 150
rect 1245 85 1338 93
rect 1109 51 1338 85
rect 1403 59 1461 147
rect 1605 117 1639 375
rect 1495 17 1529 113
rect 1579 51 1639 117
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< obsm1 >>
rect 569 320 627 329
rect 1029 320 1087 329
rect 569 292 1087 320
rect 569 283 627 292
rect 1029 283 1087 292
rect 753 184 811 193
rect 1029 184 1087 193
rect 1305 184 1363 193
rect 753 156 1363 184
rect 753 147 811 156
rect 1029 147 1087 156
rect 1305 147 1363 156
rect 845 116 903 125
rect 1397 116 1455 125
rect 845 88 1455 116
rect 845 79 903 88
rect 1397 79 1455 88
<< labels >>
rlabel locali s 1409 215 1491 265 6 A
port 1 nsew signal input
rlabel locali s 1245 199 1279 289 6 B
port 2 nsew signal input
rlabel locali s 1245 289 1361 323 6 B
port 2 nsew signal input
rlabel locali s 323 215 436 265 6 C
port 3 nsew signal input
rlabel metal1 s 0 -48 1656 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1256 21 1652 23 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 655 21 845 23 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 197 23 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 23 1652 201 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 201 1341 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1694 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1656 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 17 70 69 185 6 X
port 8 nsew signal output
rlabel locali s 17 185 66 288 6 X
port 8 nsew signal output
rlabel locali s 17 288 73 493 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1656 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 596416
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 584810
<< end >>
