magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect 4002 3832 4811 4000
rect 4041 3288 4811 3832
rect 9960 3225 10663 4000
rect 10137 2431 11093 2700
rect 10027 1997 11093 2431
<< pwell >>
rect 4208 2873 4662 3183
rect 3344 2787 4683 2873
rect 10212 1676 11018 1892
rect 10203 1590 11027 1676
<< mvnmos >>
rect 4287 3017 4407 3157
rect 4463 3017 4583 3157
rect 10291 1726 10411 1866
rect 10467 1726 10587 1866
rect 10643 1726 10763 1866
rect 10819 1726 10939 1866
<< mvpmos >>
rect 4287 3623 4407 3823
rect 4463 3623 4583 3823
rect 4287 3355 4407 3555
rect 4463 3355 4583 3555
rect 10291 2332 10411 2532
rect 10467 2332 10587 2532
rect 10643 2332 10763 2532
rect 10819 2332 10939 2532
rect 10291 2064 10411 2264
rect 10467 2064 10587 2264
rect 10643 2064 10763 2264
rect 10819 2064 10939 2264
<< mvndiff >>
rect 4234 3145 4287 3157
rect 4234 3111 4242 3145
rect 4276 3111 4287 3145
rect 4234 3077 4287 3111
rect 4234 3043 4242 3077
rect 4276 3043 4287 3077
rect 4234 3017 4287 3043
rect 4407 3145 4463 3157
rect 4407 3111 4418 3145
rect 4452 3111 4463 3145
rect 4407 3077 4463 3111
rect 4407 3043 4418 3077
rect 4452 3043 4463 3077
rect 4407 3017 4463 3043
rect 4583 3145 4636 3157
rect 4583 3111 4594 3145
rect 4628 3111 4636 3145
rect 4583 3077 4636 3111
rect 4583 3043 4594 3077
rect 4628 3043 4636 3077
rect 4583 3017 4636 3043
rect 10238 1854 10291 1866
rect 10238 1820 10246 1854
rect 10280 1820 10291 1854
rect 10238 1786 10291 1820
rect 10238 1752 10246 1786
rect 10280 1752 10291 1786
rect 10238 1726 10291 1752
rect 10411 1726 10467 1866
rect 10587 1854 10643 1866
rect 10587 1820 10598 1854
rect 10632 1820 10643 1854
rect 10587 1786 10643 1820
rect 10587 1752 10598 1786
rect 10632 1752 10643 1786
rect 10587 1726 10643 1752
rect 10763 1726 10819 1866
rect 10939 1854 10992 1866
rect 10939 1820 10950 1854
rect 10984 1820 10992 1854
rect 10939 1786 10992 1820
rect 10939 1752 10950 1786
rect 10984 1752 10992 1786
rect 10939 1726 10992 1752
<< mvpdiff >>
rect 4234 3805 4287 3823
rect 4234 3771 4242 3805
rect 4276 3771 4287 3805
rect 4234 3737 4287 3771
rect 4234 3703 4242 3737
rect 4276 3703 4287 3737
rect 4234 3669 4287 3703
rect 4234 3635 4242 3669
rect 4276 3635 4287 3669
rect 4234 3623 4287 3635
rect 4407 3805 4463 3823
rect 4407 3771 4418 3805
rect 4452 3771 4463 3805
rect 4407 3737 4463 3771
rect 4407 3703 4418 3737
rect 4452 3703 4463 3737
rect 4407 3669 4463 3703
rect 4407 3635 4418 3669
rect 4452 3635 4463 3669
rect 4407 3623 4463 3635
rect 4583 3805 4636 3823
rect 4583 3771 4594 3805
rect 4628 3771 4636 3805
rect 4583 3737 4636 3771
rect 4583 3703 4594 3737
rect 4628 3703 4636 3737
rect 4583 3669 4636 3703
rect 4583 3635 4594 3669
rect 4628 3635 4636 3669
rect 4583 3623 4636 3635
rect 4234 3543 4287 3555
rect 4234 3509 4242 3543
rect 4276 3509 4287 3543
rect 4234 3475 4287 3509
rect 4234 3441 4242 3475
rect 4276 3441 4287 3475
rect 4234 3407 4287 3441
rect 4234 3373 4242 3407
rect 4276 3373 4287 3407
rect 4234 3355 4287 3373
rect 4407 3543 4463 3555
rect 4407 3509 4418 3543
rect 4452 3509 4463 3543
rect 4407 3475 4463 3509
rect 4407 3441 4418 3475
rect 4452 3441 4463 3475
rect 4407 3407 4463 3441
rect 4407 3373 4418 3407
rect 4452 3373 4463 3407
rect 4407 3355 4463 3373
rect 4583 3543 4636 3555
rect 4583 3509 4594 3543
rect 4628 3509 4636 3543
rect 4583 3475 4636 3509
rect 4583 3441 4594 3475
rect 4628 3441 4636 3475
rect 4583 3407 4636 3441
rect 4583 3373 4594 3407
rect 4628 3373 4636 3407
rect 4583 3355 4636 3373
rect 10238 2514 10291 2532
rect 10238 2480 10246 2514
rect 10280 2480 10291 2514
rect 10238 2446 10291 2480
rect 10238 2412 10246 2446
rect 10280 2412 10291 2446
rect 10238 2378 10291 2412
rect 10238 2344 10246 2378
rect 10280 2344 10291 2378
rect 10238 2332 10291 2344
rect 10411 2514 10467 2532
rect 10411 2480 10422 2514
rect 10456 2480 10467 2514
rect 10411 2446 10467 2480
rect 10411 2412 10422 2446
rect 10456 2412 10467 2446
rect 10411 2378 10467 2412
rect 10411 2344 10422 2378
rect 10456 2344 10467 2378
rect 10411 2332 10467 2344
rect 10587 2514 10643 2532
rect 10587 2480 10598 2514
rect 10632 2480 10643 2514
rect 10587 2446 10643 2480
rect 10587 2412 10598 2446
rect 10632 2412 10643 2446
rect 10587 2378 10643 2412
rect 10587 2344 10598 2378
rect 10632 2344 10643 2378
rect 10587 2332 10643 2344
rect 10763 2514 10819 2532
rect 10763 2480 10774 2514
rect 10808 2480 10819 2514
rect 10763 2446 10819 2480
rect 10763 2412 10774 2446
rect 10808 2412 10819 2446
rect 10763 2378 10819 2412
rect 10763 2344 10774 2378
rect 10808 2344 10819 2378
rect 10763 2332 10819 2344
rect 10939 2514 10992 2532
rect 10939 2480 10950 2514
rect 10984 2480 10992 2514
rect 10939 2446 10992 2480
rect 10939 2412 10950 2446
rect 10984 2412 10992 2446
rect 10939 2378 10992 2412
rect 10939 2344 10950 2378
rect 10984 2344 10992 2378
rect 10939 2332 10992 2344
rect 10238 2252 10291 2264
rect 10238 2218 10246 2252
rect 10280 2218 10291 2252
rect 10238 2184 10291 2218
rect 10238 2150 10246 2184
rect 10280 2150 10291 2184
rect 10238 2116 10291 2150
rect 10238 2082 10246 2116
rect 10280 2082 10291 2116
rect 10238 2064 10291 2082
rect 10411 2252 10467 2264
rect 10411 2218 10422 2252
rect 10456 2218 10467 2252
rect 10411 2184 10467 2218
rect 10411 2150 10422 2184
rect 10456 2150 10467 2184
rect 10411 2116 10467 2150
rect 10411 2082 10422 2116
rect 10456 2082 10467 2116
rect 10411 2064 10467 2082
rect 10587 2252 10643 2264
rect 10587 2218 10598 2252
rect 10632 2218 10643 2252
rect 10587 2184 10643 2218
rect 10587 2150 10598 2184
rect 10632 2150 10643 2184
rect 10587 2116 10643 2150
rect 10587 2082 10598 2116
rect 10632 2082 10643 2116
rect 10587 2064 10643 2082
rect 10763 2252 10819 2264
rect 10763 2218 10774 2252
rect 10808 2218 10819 2252
rect 10763 2184 10819 2218
rect 10763 2150 10774 2184
rect 10808 2150 10819 2184
rect 10763 2116 10819 2150
rect 10763 2082 10774 2116
rect 10808 2082 10819 2116
rect 10763 2064 10819 2082
rect 10939 2252 10992 2264
rect 10939 2218 10950 2252
rect 10984 2218 10992 2252
rect 10939 2184 10992 2218
rect 10939 2150 10950 2184
rect 10984 2150 10992 2184
rect 10939 2116 10992 2150
rect 10939 2082 10950 2116
rect 10984 2082 10992 2116
rect 10939 2064 10992 2082
<< mvndiffc >>
rect 4242 3111 4276 3145
rect 4242 3043 4276 3077
rect 4418 3111 4452 3145
rect 4418 3043 4452 3077
rect 4594 3111 4628 3145
rect 4594 3043 4628 3077
rect 10246 1820 10280 1854
rect 10246 1752 10280 1786
rect 10598 1820 10632 1854
rect 10598 1752 10632 1786
rect 10950 1820 10984 1854
rect 10950 1752 10984 1786
<< mvpdiffc >>
rect 4242 3771 4276 3805
rect 4242 3703 4276 3737
rect 4242 3635 4276 3669
rect 4418 3771 4452 3805
rect 4418 3703 4452 3737
rect 4418 3635 4452 3669
rect 4594 3771 4628 3805
rect 4594 3703 4628 3737
rect 4594 3635 4628 3669
rect 4242 3509 4276 3543
rect 4242 3441 4276 3475
rect 4242 3373 4276 3407
rect 4418 3509 4452 3543
rect 4418 3441 4452 3475
rect 4418 3373 4452 3407
rect 4594 3509 4628 3543
rect 4594 3441 4628 3475
rect 4594 3373 4628 3407
rect 10246 2480 10280 2514
rect 10246 2412 10280 2446
rect 10246 2344 10280 2378
rect 10422 2480 10456 2514
rect 10422 2412 10456 2446
rect 10422 2344 10456 2378
rect 10598 2480 10632 2514
rect 10598 2412 10632 2446
rect 10598 2344 10632 2378
rect 10774 2480 10808 2514
rect 10774 2412 10808 2446
rect 10774 2344 10808 2378
rect 10950 2480 10984 2514
rect 10950 2412 10984 2446
rect 10950 2344 10984 2378
rect 10246 2218 10280 2252
rect 10246 2150 10280 2184
rect 10246 2082 10280 2116
rect 10422 2218 10456 2252
rect 10422 2150 10456 2184
rect 10422 2082 10456 2116
rect 10598 2218 10632 2252
rect 10598 2150 10632 2184
rect 10598 2082 10632 2116
rect 10774 2218 10808 2252
rect 10774 2150 10808 2184
rect 10774 2082 10808 2116
rect 10950 2218 10984 2252
rect 10950 2150 10984 2184
rect 10950 2082 10984 2116
<< mvpsubdiff >>
rect 3370 2813 3394 2847
rect 3428 2813 3465 2847
rect 3499 2813 3536 2847
rect 3570 2813 3607 2847
rect 3641 2813 3678 2847
rect 3712 2813 3749 2847
rect 3783 2813 3820 2847
rect 3854 2813 3891 2847
rect 3925 2813 3962 2847
rect 3996 2813 4033 2847
rect 4067 2813 4104 2847
rect 4138 2813 4175 2847
rect 4209 2813 4246 2847
rect 4280 2813 4317 2847
rect 4351 2813 4388 2847
rect 4422 2813 4459 2847
rect 4493 2813 4529 2847
rect 4563 2813 4599 2847
rect 4633 2813 4657 2847
rect 10229 1616 10253 1650
rect 10287 1616 10322 1650
rect 10356 1616 10391 1650
rect 10425 1616 10460 1650
rect 10494 1616 10529 1650
rect 10563 1616 10598 1650
rect 10632 1616 10667 1650
rect 10701 1616 10736 1650
rect 10770 1616 10805 1650
rect 10839 1616 10874 1650
rect 10908 1616 10943 1650
rect 10977 1616 11001 1650
<< mvnsubdiff >>
rect 4069 3899 4103 3933
rect 4137 3899 4171 3933
rect 4205 3899 4239 3933
rect 4273 3899 4307 3933
rect 4341 3899 4375 3933
rect 4409 3899 4443 3933
rect 4477 3899 4511 3933
rect 4545 3899 4579 3933
rect 4613 3899 4647 3933
rect 4681 3899 4744 3933
rect 10203 2600 10227 2634
rect 10261 2600 10302 2634
rect 10336 2600 10377 2634
rect 10411 2600 10451 2634
rect 10485 2600 10525 2634
rect 10559 2600 10599 2634
rect 10633 2600 10673 2634
rect 10707 2600 10747 2634
rect 10781 2600 10821 2634
rect 10855 2600 10895 2634
rect 10929 2600 10969 2634
rect 11003 2600 11027 2634
<< mvpsubdiffcont >>
rect 3394 2813 3428 2847
rect 3465 2813 3499 2847
rect 3536 2813 3570 2847
rect 3607 2813 3641 2847
rect 3678 2813 3712 2847
rect 3749 2813 3783 2847
rect 3820 2813 3854 2847
rect 3891 2813 3925 2847
rect 3962 2813 3996 2847
rect 4033 2813 4067 2847
rect 4104 2813 4138 2847
rect 4175 2813 4209 2847
rect 4246 2813 4280 2847
rect 4317 2813 4351 2847
rect 4388 2813 4422 2847
rect 4459 2813 4493 2847
rect 4529 2813 4563 2847
rect 4599 2813 4633 2847
rect 10253 1616 10287 1650
rect 10322 1616 10356 1650
rect 10391 1616 10425 1650
rect 10460 1616 10494 1650
rect 10529 1616 10563 1650
rect 10598 1616 10632 1650
rect 10667 1616 10701 1650
rect 10736 1616 10770 1650
rect 10805 1616 10839 1650
rect 10874 1616 10908 1650
rect 10943 1616 10977 1650
<< mvnsubdiffcont >>
rect 4103 3899 4137 3933
rect 4171 3899 4205 3933
rect 4239 3899 4273 3933
rect 4307 3899 4341 3933
rect 4375 3899 4409 3933
rect 4443 3899 4477 3933
rect 4511 3899 4545 3933
rect 4579 3899 4613 3933
rect 4647 3899 4681 3933
rect 10227 2600 10261 2634
rect 10302 2600 10336 2634
rect 10377 2600 10411 2634
rect 10451 2600 10485 2634
rect 10525 2600 10559 2634
rect 10599 2600 10633 2634
rect 10673 2600 10707 2634
rect 10747 2600 10781 2634
rect 10821 2600 10855 2634
rect 10895 2600 10929 2634
rect 10969 2600 11003 2634
<< poly >>
rect 4287 3823 4407 3849
rect 4463 3823 4583 3849
rect 4287 3555 4407 3623
rect 4463 3555 4583 3623
rect 4287 3307 4407 3355
rect 4287 3273 4329 3307
rect 4363 3273 4407 3307
rect 4287 3239 4407 3273
rect 4287 3205 4329 3239
rect 4363 3205 4407 3239
rect 4287 3157 4407 3205
rect 4463 3307 4583 3355
rect 4463 3273 4507 3307
rect 4541 3273 4583 3307
rect 4463 3239 4583 3273
rect 4463 3205 4507 3239
rect 4541 3205 4583 3239
rect 4463 3157 4583 3205
rect 4287 2991 4407 3017
rect 4463 2991 4583 3017
rect 10291 2532 10411 2558
rect 10467 2532 10587 2558
rect 10643 2532 10763 2558
rect 10819 2532 10939 2558
rect 10291 2264 10411 2332
rect 10467 2264 10587 2332
rect 10643 2264 10763 2332
rect 10819 2264 10939 2332
rect 10291 2016 10411 2064
rect 10291 1982 10336 2016
rect 10370 1982 10411 2016
rect 10291 1948 10411 1982
rect 10291 1914 10336 1948
rect 10370 1914 10411 1948
rect 10291 1866 10411 1914
rect 10467 2016 10587 2064
rect 10467 1982 10507 2016
rect 10541 1982 10587 2016
rect 10467 1948 10587 1982
rect 10467 1914 10507 1948
rect 10541 1914 10587 1948
rect 10467 1866 10587 1914
rect 10643 2016 10763 2064
rect 10643 1982 10689 2016
rect 10723 1982 10763 2016
rect 10643 1948 10763 1982
rect 10643 1914 10689 1948
rect 10723 1914 10763 1948
rect 10643 1866 10763 1914
rect 10819 2016 10939 2064
rect 10819 1982 10860 2016
rect 10894 1982 10939 2016
rect 10819 1948 10939 1982
rect 10819 1914 10860 1948
rect 10894 1914 10939 1948
rect 10819 1866 10939 1914
rect 10291 1700 10411 1726
rect 10467 1700 10587 1726
rect 10643 1700 10763 1726
rect 10819 1700 10939 1726
<< polycont >>
rect 4329 3273 4363 3307
rect 4329 3205 4363 3239
rect 4507 3273 4541 3307
rect 4507 3205 4541 3239
rect 10336 1982 10370 2016
rect 10336 1914 10370 1948
rect 10507 1982 10541 2016
rect 10507 1914 10541 1948
rect 10689 1982 10723 2016
rect 10689 1914 10723 1948
rect 10860 1982 10894 2016
rect 10860 1914 10894 1948
<< locali >>
rect 4069 3899 4084 3933
rect 4137 3899 4161 3933
rect 4205 3899 4238 3933
rect 4273 3899 4307 3933
rect 4349 3899 4375 3933
rect 4426 3899 4443 3933
rect 4503 3899 4511 3933
rect 4545 3899 4546 3933
rect 4613 3899 4622 3933
rect 4681 3899 4698 3933
rect 4732 3899 4744 3933
rect 4242 3805 4276 3823
rect 4242 3737 4276 3771
rect 4242 3669 4276 3703
rect 4242 3543 4276 3635
rect 4242 3475 4276 3509
rect 4242 3407 4276 3441
rect 4242 3314 4276 3373
rect 4418 3805 4452 3817
rect 4418 3737 4452 3745
rect 4418 3669 4452 3703
rect 4418 3543 4452 3635
rect 4418 3475 4452 3509
rect 4418 3407 4452 3441
rect 4418 3357 4452 3373
rect 4594 3805 4628 3823
rect 4594 3737 4628 3771
rect 4594 3669 4628 3703
rect 4594 3543 4628 3635
rect 4594 3475 4628 3509
rect 4594 3407 4628 3441
rect 4594 3314 4628 3373
rect 4270 3280 4276 3314
rect 4236 3242 4276 3280
rect 4270 3208 4276 3242
rect 4242 3145 4276 3208
rect 4313 3273 4329 3307
rect 4370 3280 4379 3307
rect 4363 3273 4379 3280
rect 4313 3242 4379 3273
rect 4313 3239 4336 3242
rect 4313 3205 4329 3239
rect 4370 3208 4379 3242
rect 4363 3205 4379 3208
rect 4491 3280 4492 3307
rect 4491 3273 4507 3280
rect 4541 3273 4557 3307
rect 4491 3242 4557 3273
rect 4491 3208 4492 3242
rect 4526 3239 4557 3242
rect 4491 3205 4507 3208
rect 4541 3205 4557 3239
rect 4594 3242 4628 3280
rect 4242 3077 4276 3111
rect 4242 3027 4276 3043
rect 4418 3145 4452 3161
rect 4418 3100 4452 3111
rect 4418 3028 4452 3043
rect 4594 3145 4628 3208
rect 4594 3077 4628 3111
rect 4594 3027 4628 3043
rect 3370 2813 3394 2847
rect 3428 2813 3464 2847
rect 3499 2813 3536 2847
rect 3575 2813 3607 2847
rect 3652 2813 3678 2847
rect 3729 2813 3749 2847
rect 3806 2813 3820 2847
rect 3883 2813 3891 2847
rect 3925 2813 3926 2847
rect 3960 2813 3962 2847
rect 3996 2813 4003 2847
rect 4067 2813 4079 2847
rect 4138 2813 4155 2847
rect 4209 2813 4231 2847
rect 4280 2813 4307 2847
rect 4351 2813 4383 2847
rect 4422 2813 4459 2847
rect 4493 2813 4529 2847
rect 4569 2813 4599 2847
rect 4645 2813 4657 2847
rect 10203 2600 10215 2634
rect 10261 2600 10292 2634
rect 10336 2600 10369 2634
rect 10411 2600 10446 2634
rect 10485 2600 10523 2634
rect 10559 2600 10599 2634
rect 10634 2600 10673 2634
rect 10711 2600 10747 2634
rect 10787 2600 10821 2634
rect 10863 2600 10895 2634
rect 10939 2600 10969 2634
rect 11015 2600 11027 2634
rect 10246 2514 10280 2526
rect 10246 2446 10280 2454
rect 10246 2378 10280 2412
rect 10246 2252 10280 2344
rect 10246 2184 10280 2218
rect 10246 2116 10280 2150
rect 10246 2066 10280 2082
rect 10422 2514 10456 2532
rect 10422 2446 10456 2480
rect 10422 2378 10456 2412
rect 10422 2252 10456 2344
rect 10422 2184 10456 2218
rect 10422 2116 10456 2150
rect 10320 1982 10336 1986
rect 10370 1982 10386 2016
rect 10320 1948 10386 1982
rect 10370 1914 10386 1948
rect 10422 1967 10456 2082
rect 10598 2514 10632 2526
rect 10598 2446 10632 2454
rect 10598 2378 10632 2412
rect 10598 2252 10632 2344
rect 10598 2184 10632 2218
rect 10598 2116 10632 2150
rect 10598 2066 10632 2082
rect 10774 2514 10808 2532
rect 10774 2446 10808 2480
rect 10774 2378 10808 2412
rect 10774 2252 10808 2344
rect 10774 2184 10808 2218
rect 10774 2116 10808 2121
rect 10950 2514 10984 2526
rect 10950 2446 10984 2454
rect 10950 2378 10984 2412
rect 10950 2252 10984 2344
rect 10950 2184 10984 2218
rect 10950 2116 10984 2150
rect 10950 2066 10984 2082
rect 10422 1895 10456 1933
rect 10491 1982 10507 2016
rect 10541 1982 10689 2016
rect 10723 1982 10739 2016
rect 10491 1969 10739 1982
rect 10491 1948 10521 1969
rect 10491 1914 10507 1948
rect 10555 1935 10593 1969
rect 10627 1948 10739 1969
rect 10627 1935 10689 1948
rect 10541 1914 10689 1935
rect 10723 1914 10739 1948
rect 10246 1854 10280 1870
rect 10422 1843 10456 1861
rect 10280 1820 10456 1843
rect 10246 1809 10456 1820
rect 10598 1854 10632 1870
rect 10598 1809 10632 1820
rect 10774 1843 10808 2049
rect 10844 2003 10860 2016
rect 10894 2003 10910 2016
rect 10894 1982 10916 2003
rect 10878 1969 10916 1982
rect 10844 1948 10910 1969
rect 10844 1914 10860 1948
rect 10894 1914 10910 1948
rect 10950 1854 10984 1870
rect 10774 1820 10950 1843
rect 10774 1809 10984 1820
rect 10246 1786 10285 1809
rect 10280 1752 10285 1786
rect 10246 1736 10285 1752
rect 10598 1737 10632 1752
rect 10945 1786 10984 1809
rect 10945 1752 10950 1786
rect 10945 1736 10984 1752
rect 10229 1616 10241 1650
rect 10287 1616 10315 1650
rect 10356 1616 10389 1650
rect 10425 1616 10460 1650
rect 10497 1616 10529 1650
rect 10571 1616 10598 1650
rect 10645 1616 10667 1650
rect 10719 1616 10736 1650
rect 10793 1616 10805 1650
rect 10867 1616 10874 1650
rect 10941 1616 10943 1650
rect 10977 1616 10981 1650
<< viali >>
rect 4084 3899 4103 3933
rect 4103 3899 4118 3933
rect 4161 3899 4171 3933
rect 4171 3899 4195 3933
rect 4238 3899 4239 3933
rect 4239 3899 4272 3933
rect 4315 3899 4341 3933
rect 4341 3899 4349 3933
rect 4392 3899 4409 3933
rect 4409 3899 4426 3933
rect 4469 3899 4477 3933
rect 4477 3899 4503 3933
rect 4546 3899 4579 3933
rect 4579 3899 4580 3933
rect 4622 3899 4647 3933
rect 4647 3899 4656 3933
rect 4698 3899 4732 3933
rect 4418 3817 4452 3851
rect 4418 3771 4452 3779
rect 4418 3745 4452 3771
rect 4236 3280 4270 3314
rect 4336 3307 4370 3314
rect 4492 3307 4526 3314
rect 4236 3208 4270 3242
rect 4336 3280 4363 3307
rect 4363 3280 4370 3307
rect 4336 3239 4370 3242
rect 4336 3208 4363 3239
rect 4363 3208 4370 3239
rect 4492 3280 4507 3307
rect 4507 3280 4526 3307
rect 4492 3239 4526 3242
rect 4492 3208 4507 3239
rect 4507 3208 4526 3239
rect 4594 3280 4628 3314
rect 4594 3208 4628 3242
rect 4418 3077 4452 3100
rect 4418 3066 4452 3077
rect 4418 2994 4452 3028
rect 3464 2813 3465 2847
rect 3465 2813 3498 2847
rect 3541 2813 3570 2847
rect 3570 2813 3575 2847
rect 3618 2813 3641 2847
rect 3641 2813 3652 2847
rect 3695 2813 3712 2847
rect 3712 2813 3729 2847
rect 3772 2813 3783 2847
rect 3783 2813 3806 2847
rect 3849 2813 3854 2847
rect 3854 2813 3883 2847
rect 3926 2813 3960 2847
rect 4003 2813 4033 2847
rect 4033 2813 4037 2847
rect 4079 2813 4104 2847
rect 4104 2813 4113 2847
rect 4155 2813 4175 2847
rect 4175 2813 4189 2847
rect 4231 2813 4246 2847
rect 4246 2813 4265 2847
rect 4307 2813 4317 2847
rect 4317 2813 4341 2847
rect 4383 2813 4388 2847
rect 4388 2813 4417 2847
rect 4459 2813 4493 2847
rect 4535 2813 4563 2847
rect 4563 2813 4569 2847
rect 4611 2813 4633 2847
rect 4633 2813 4645 2847
rect 10215 2600 10227 2634
rect 10227 2600 10249 2634
rect 10292 2600 10302 2634
rect 10302 2600 10326 2634
rect 10369 2600 10377 2634
rect 10377 2600 10403 2634
rect 10446 2600 10451 2634
rect 10451 2600 10480 2634
rect 10523 2600 10525 2634
rect 10525 2600 10557 2634
rect 10600 2600 10633 2634
rect 10633 2600 10634 2634
rect 10677 2600 10707 2634
rect 10707 2600 10711 2634
rect 10753 2600 10781 2634
rect 10781 2600 10787 2634
rect 10829 2600 10855 2634
rect 10855 2600 10863 2634
rect 10905 2600 10929 2634
rect 10929 2600 10939 2634
rect 10981 2600 11003 2634
rect 11003 2600 11015 2634
rect 10246 2526 10280 2560
rect 10246 2480 10280 2488
rect 10246 2454 10280 2480
rect 10320 2016 10354 2020
rect 10320 1986 10336 2016
rect 10336 1986 10354 2016
rect 10320 1914 10336 1948
rect 10336 1914 10354 1948
rect 10598 2526 10632 2560
rect 10598 2480 10632 2488
rect 10598 2454 10632 2480
rect 10774 2150 10808 2155
rect 10774 2121 10808 2150
rect 10774 2082 10808 2083
rect 10774 2049 10808 2082
rect 10950 2526 10984 2560
rect 10950 2480 10984 2488
rect 10950 2454 10984 2480
rect 10422 1933 10456 1967
rect 10521 1948 10555 1969
rect 10521 1935 10541 1948
rect 10541 1935 10555 1948
rect 10593 1935 10627 1969
rect 10422 1861 10456 1895
rect 10844 1982 10860 2003
rect 10860 1982 10878 2003
rect 10844 1969 10878 1982
rect 10916 1969 10950 2003
rect 10598 1786 10632 1809
rect 10598 1775 10632 1786
rect 10598 1703 10632 1737
rect 10241 1616 10253 1650
rect 10253 1616 10275 1650
rect 10315 1616 10322 1650
rect 10322 1616 10349 1650
rect 10389 1616 10391 1650
rect 10391 1616 10423 1650
rect 10463 1616 10494 1650
rect 10494 1616 10497 1650
rect 10537 1616 10563 1650
rect 10563 1616 10571 1650
rect 10611 1616 10632 1650
rect 10632 1616 10645 1650
rect 10685 1616 10701 1650
rect 10701 1616 10719 1650
rect 10759 1616 10770 1650
rect 10770 1616 10793 1650
rect 10833 1616 10839 1650
rect 10839 1616 10867 1650
rect 10907 1616 10908 1650
rect 10908 1616 10941 1650
rect 10981 1616 11015 1650
<< metal1 >>
rect 68 3933 4839 4000
rect 68 3899 4084 3933
rect 4118 3899 4161 3933
rect 4195 3899 4238 3933
rect 4272 3899 4315 3933
rect 4349 3899 4392 3933
rect 4426 3899 4469 3933
rect 4503 3899 4546 3933
rect 4580 3899 4622 3933
rect 4656 3899 4698 3933
rect 4732 3899 4839 3933
rect 68 3851 4839 3899
rect 68 3817 4418 3851
rect 4452 3817 4839 3851
rect 68 3779 4839 3817
rect 10001 3801 10740 4000
rect 68 3745 4418 3779
rect 4452 3745 4839 3779
tri 10009 3767 10043 3801 nw
tri 10169 3767 10203 3801 ne
tri 10465 3767 10499 3801 nw
tri 10629 3767 10663 3801 ne
tri 10696 3767 10730 3801 ne
rect 11495 3762 12100 3985
rect 68 3732 4839 3745
rect 4227 3320 4279 3326
rect 4227 3254 4279 3268
rect 4227 3196 4279 3202
rect 4327 3320 4379 3326
rect 4327 3254 4379 3268
rect 4327 3196 4379 3202
rect 4483 3320 4535 3326
rect 4483 3254 4535 3268
rect 4483 3196 4535 3202
rect 4585 3320 4637 3326
rect 4585 3254 4637 3268
rect 4585 3196 4637 3202
tri 10069 3223 10075 3229 se
tri 10593 3225 10597 3229 sw
rect 10069 3217 10121 3223
rect 10069 3153 10121 3165
rect 3951 3106 4683 3112
rect 3951 3054 4106 3106
rect 4158 3100 4683 3106
rect 4158 3066 4418 3100
rect 4452 3066 4683 3100
rect 10069 3095 10121 3101
rect 10149 3219 10201 3225
rect 10149 3153 10201 3167
rect 10149 3095 10201 3101
rect 10467 3219 10519 3225
rect 10593 3223 10597 3225
tri 10597 3223 10599 3225 sw
rect 10467 3153 10519 3167
rect 10467 3095 10519 3101
rect 10547 3217 10599 3223
rect 10547 3153 10599 3165
rect 10547 3095 10599 3101
tri 10069 3089 10075 3095 ne
tri 10593 3089 10599 3095 nw
rect 4158 3054 4683 3066
rect 3951 3031 4683 3054
rect 3951 2979 4106 3031
rect 4158 3028 4683 3031
rect 4158 2994 4418 3028
rect 4452 2994 4683 3028
rect 4158 2979 4683 2994
rect 3951 2955 4683 2979
rect 3951 2903 4106 2955
rect 4158 2903 4683 2955
rect 3452 2897 4683 2903
tri 3362 2847 3412 2897 ne
rect 3412 2847 4683 2897
rect 10358 3053 10437 3059
rect 10358 3001 10371 3053
rect 10423 3001 10437 3053
rect 10358 2987 10437 3001
rect 10358 2935 10371 2987
rect 10423 2935 10437 2987
rect 10358 2921 10437 2935
rect 10358 2869 10371 2921
rect 10423 2869 10437 2921
rect 10358 2863 10437 2869
tri 3412 2835 3424 2847 ne
rect 3424 2835 3464 2847
tri 3424 2813 3446 2835 ne
rect 3446 2813 3464 2835
rect 3498 2813 3541 2847
rect 3575 2813 3618 2847
rect 3652 2813 3695 2847
rect 3729 2813 3772 2847
rect 3806 2813 3849 2847
rect 3883 2813 3926 2847
rect 3960 2813 4003 2847
rect 4037 2813 4079 2847
rect 4113 2813 4155 2847
rect 4189 2813 4231 2847
rect 4265 2813 4307 2847
rect 4341 2813 4383 2847
rect 4417 2813 4459 2847
rect 4493 2813 4535 2847
rect 4569 2813 4611 2847
rect 4645 2813 4683 2847
tri 3446 2807 3452 2813 ne
rect 3452 2807 4683 2813
rect 10467 2829 12109 2835
tri 10039 2731 10091 2783 se
rect 10091 2731 10208 2783
rect 10260 2731 10272 2783
rect 10324 2731 10330 2783
rect 10519 2783 12109 2829
rect 12161 2783 12173 2835
rect 12225 2783 12231 2835
rect 10467 2765 10519 2777
tri 10003 2695 10039 2731 se
rect 10039 2707 10089 2731
tri 10089 2707 10113 2731 nw
tri 10519 2749 10553 2783 nw
rect 10467 2707 10519 2713
tri 11018 2707 11024 2713 se
rect 10039 2695 10077 2707
tri 10077 2695 10089 2707 nw
tri 11006 2695 11018 2707 se
rect 11018 2695 11024 2707
tri 9985 2677 10003 2695 se
rect 10003 2677 10016 2695
rect 99 2628 266 2672
rect 4327 2625 4333 2677
rect 4385 2625 4397 2677
rect 4449 2625 4455 2677
tri 9981 2673 9985 2677 se
rect 9985 2673 10016 2677
rect 9846 2634 10016 2673
tri 10016 2634 10077 2695 nw
tri 10955 2644 11006 2695 se
rect 11006 2644 11024 2695
rect 10203 2634 11027 2644
rect 9846 2621 10003 2634
tri 10003 2621 10016 2634 nw
rect 10203 2600 10215 2634
rect 10249 2600 10292 2634
rect 10326 2600 10369 2634
rect 10403 2600 10446 2634
rect 10480 2600 10523 2634
rect 10557 2600 10600 2634
rect 10634 2600 10677 2634
rect 10711 2600 10753 2634
rect 10787 2600 10829 2634
rect 10863 2600 10905 2634
rect 10939 2600 10981 2634
rect 11015 2600 11027 2634
rect 91 2545 4489 2597
rect 4541 2545 4553 2597
rect 4605 2545 4799 2597
rect 10203 2560 11027 2600
rect 10203 2526 10246 2560
rect 10280 2526 10598 2560
rect 10632 2526 10950 2560
rect 10984 2526 11027 2560
rect 4227 2465 4233 2517
rect 4285 2465 4297 2517
rect 4349 2465 4799 2517
rect 8334 2501 10021 2507
rect 8386 2488 10021 2501
tri 10021 2488 10040 2507 sw
rect 10203 2488 11027 2526
rect 8386 2462 10040 2488
tri 10040 2462 10066 2488 sw
rect 8386 2455 10066 2462
rect 8386 2454 8419 2455
tri 8419 2454 8420 2455 nw
tri 9999 2454 10000 2455 ne
rect 10000 2454 10066 2455
tri 10066 2454 10074 2462 sw
rect 10203 2454 10246 2488
rect 10280 2454 10598 2488
rect 10632 2454 10950 2488
rect 10984 2454 11027 2488
rect 8334 2437 8386 2449
rect 397 2393 483 2427
tri 8386 2421 8419 2454 nw
tri 10000 2421 10033 2454 ne
rect 10033 2421 10074 2454
tri 10033 2388 10066 2421 ne
rect 10066 2388 10074 2421
tri 10074 2388 10140 2454 sw
rect 10203 2441 11027 2454
rect 8334 2379 8386 2385
tri 10066 2379 10075 2388 ne
rect 10075 2379 10140 2388
tri 10075 2366 10088 2379 ne
rect 10088 2167 10140 2379
tri 10930 2347 11024 2441 ne
rect 11285 2355 11293 2357
tri 11293 2355 11295 2357 nw
rect 11024 2347 11285 2355
tri 11285 2347 11293 2355 nw
rect 10278 2323 10330 2329
rect 11402 2323 11454 2329
rect 10278 2259 10330 2271
tri 10330 2253 10364 2287 sw
tri 11368 2253 11402 2287 se
rect 11402 2259 11454 2271
rect 10330 2207 11402 2253
rect 10278 2201 11454 2207
tri 10140 2167 10162 2189 sw
tri 10088 2155 10100 2167 ne
rect 10100 2155 10162 2167
tri 10162 2155 10174 2167 sw
rect 10768 2155 10814 2167
tri 10100 2139 10116 2155 ne
rect 10116 2139 10174 2155
tri 10174 2139 10190 2155 sw
tri 10116 2121 10134 2139 ne
rect 10134 2121 10598 2139
tri 10598 2121 10616 2139 sw
rect 10768 2121 10774 2155
rect 10808 2121 10814 2155
tri 10134 2115 10140 2121 ne
rect 10140 2115 10616 2121
tri 10140 2104 10151 2115 ne
rect 10151 2104 10616 2115
rect 265 2069 398 2104
tri 10151 2087 10168 2104 ne
rect 10168 2087 10616 2104
tri 10616 2087 10650 2121 sw
rect 10768 2089 10814 2121
tri 10814 2089 10848 2123 sw
tri 10576 2083 10580 2087 ne
rect 10580 2083 10650 2087
tri 10650 2083 10654 2087 sw
rect 10768 2083 12041 2089
tri 10580 2069 10594 2083 ne
rect 10594 2069 10654 2083
tri 10594 2049 10614 2069 ne
rect 10614 2049 10654 2069
tri 10654 2049 10688 2083 sw
rect 10768 2049 10774 2083
rect 10808 2049 12041 2083
tri 10614 2032 10631 2049 ne
rect 10631 2032 10688 2049
rect 10003 2026 10360 2032
rect 10055 2020 10360 2026
rect 10055 1994 10320 2020
rect 10055 1986 10081 1994
tri 10081 1986 10089 1994 nw
tri 10280 1986 10288 1994 ne
rect 10288 1986 10320 1994
rect 10354 1986 10360 2020
tri 10631 2013 10650 2032 ne
rect 10650 2031 10688 2032
tri 10688 2031 10706 2049 sw
rect 10768 2037 12041 2049
rect 10650 2013 10706 2031
tri 10706 2013 10724 2031 sw
tri 10650 2003 10660 2013 ne
rect 10660 2009 10724 2013
tri 10724 2009 10728 2013 sw
rect 10660 2003 10962 2009
rect 10055 1974 10064 1986
rect 10003 1969 10064 1974
tri 10064 1969 10081 1986 nw
tri 10288 1969 10305 1986 ne
rect 10305 1969 10360 1986
tri 10660 1979 10684 2003 ne
rect 10684 1979 10844 2003
rect 10003 1967 10062 1969
tri 10062 1967 10064 1969 nw
tri 10305 1967 10307 1969 ne
rect 10307 1967 10360 1969
rect 10003 1962 10055 1967
tri 10055 1960 10062 1967 nw
tri 10307 1960 10314 1967 ne
rect 10003 1904 10055 1910
rect 10314 1948 10360 1967
rect 10314 1914 10320 1948
rect 10354 1914 10360 1948
rect 10314 1902 10360 1914
rect 10416 1967 10462 1979
tri 10684 1975 10688 1979 ne
rect 10688 1975 10844 1979
rect 10416 1933 10422 1967
rect 10456 1933 10462 1967
rect 10509 1969 10639 1975
tri 10688 1969 10694 1975 ne
rect 10694 1969 10844 1975
rect 10878 1969 10916 2003
rect 10950 1969 10962 2003
rect 10509 1935 10521 1969
rect 10555 1935 10593 1969
rect 10627 1935 10639 1969
tri 10694 1957 10706 1969 ne
rect 10706 1957 10962 1969
rect 12230 1946 12377 1995
rect 10416 1929 10462 1933
tri 10462 1929 10468 1935 sw
rect 10509 1929 10639 1935
rect 10416 1901 10468 1929
tri 10468 1901 10496 1929 sw
rect 10416 1895 11423 1901
rect 8334 1875 8386 1881
tri 8308 1809 8334 1835 se
rect 10416 1861 10422 1895
rect 10456 1861 11423 1895
rect 10416 1849 11423 1861
rect 8334 1811 8386 1823
tri 11368 1821 11396 1849 ne
rect 11396 1821 11402 1849
tri 8300 1801 8308 1809 se
rect 8308 1801 8334 1809
rect 7558 1759 8334 1801
tri 7536 1737 7558 1759 se
rect 7558 1753 8386 1759
rect 10203 1815 11027 1821
tri 11396 1815 11402 1821 ne
rect 10203 1763 10371 1815
rect 10423 1809 11027 1815
rect 10423 1775 10598 1809
rect 10632 1775 11027 1809
rect 10423 1763 11027 1775
rect 7558 1737 7628 1753
tri 7628 1737 7644 1753 nw
rect 10203 1740 11027 1763
tri 7524 1725 7536 1737 se
rect 7536 1725 7616 1737
tri 7616 1725 7628 1737 nw
rect 6686 1673 6692 1725
rect 6744 1673 6756 1725
rect 6808 1673 7610 1725
tri 7610 1719 7616 1725 nw
rect 8233 1673 8665 1725
rect 10203 1688 10371 1740
rect 10423 1737 11027 1740
rect 10423 1703 10598 1737
rect 10632 1703 11027 1737
rect 10423 1688 11027 1703
rect 10203 1664 11027 1688
rect 10203 1650 10371 1664
rect 10423 1650 11027 1664
rect 8232 1593 8421 1645
rect 9465 1593 9471 1645
rect 9523 1593 9535 1645
rect 9587 1593 9593 1645
rect 10203 1616 10241 1650
rect 10275 1616 10315 1650
rect 10349 1616 10371 1650
rect 10423 1616 10463 1650
rect 10497 1616 10537 1650
rect 10571 1616 10611 1650
rect 10645 1616 10685 1650
rect 10719 1616 10759 1650
rect 10793 1616 10833 1650
rect 10867 1616 10907 1650
rect 10941 1616 10981 1650
rect 11015 1616 11027 1650
rect 10203 1612 10371 1616
rect 10423 1612 11027 1616
rect 10203 1606 11027 1612
tri 7629 1525 7667 1563 se
rect 7667 1525 9933 1563
tri 7615 1511 7629 1525 se
rect 7629 1511 7709 1525
tri 7709 1511 7723 1525 nw
tri 9913 1511 9927 1525 ne
rect 9927 1511 9933 1525
rect 9985 1511 9997 1563
rect 10049 1511 10055 1563
rect 10186 1513 10192 1565
rect 10244 1513 10256 1565
rect 10308 1513 10853 1565
tri 7601 1497 7615 1511 se
rect 7615 1497 7695 1511
tri 7695 1497 7709 1511 nw
rect 4726 1491 5712 1497
rect 4778 1445 5712 1491
rect 7520 1479 7677 1497
tri 7677 1479 7695 1497 nw
rect 6894 1468 6906 1479
rect 7520 1477 7675 1479
tri 7675 1477 7677 1479 nw
rect 7520 1468 7666 1477
tri 7666 1468 7675 1477 nw
rect 7520 1452 7650 1468
tri 7650 1452 7666 1468 nw
rect 9158 1452 9175 1477
rect 7520 1445 7643 1452
tri 7643 1445 7650 1452 nw
rect 4778 1439 4784 1445
rect 4726 1427 4784 1439
rect 265 1382 375 1423
rect 4778 1417 4784 1427
tri 4784 1417 4812 1445 nw
tri 4778 1411 4784 1417 nw
rect 4726 1369 4778 1375
rect 5706 1365 5712 1417
rect 5764 1365 5776 1417
rect 5828 1365 5834 1417
rect 8255 1365 10855 1417
rect 288 1322 9419 1337
tri 9419 1322 9434 1337 sw
rect 288 1285 9434 1322
tri 9434 1285 9471 1322 sw
tri 9397 1270 9412 1285 ne
rect 9412 1270 9471 1285
tri 9471 1270 9486 1285 sw
rect 9541 1270 9547 1322
rect 9599 1270 9611 1322
rect 9663 1270 11102 1322
rect 11154 1270 11166 1322
rect 11218 1270 11224 1322
tri 9412 1211 9471 1270 ne
rect 9471 1241 9486 1270
tri 9486 1241 9515 1270 sw
rect 9471 1211 9635 1241
tri 9471 1189 9493 1211 ne
rect 9493 1189 9635 1211
rect 10938 793 10969 804
rect 12738 793 12783 797
rect 4040 189 4149 195
rect 4040 137 4069 189
rect 4121 137 4149 189
rect 4040 124 4149 137
rect 4040 72 4069 124
rect 4121 72 4149 124
rect 4040 58 4149 72
rect 1179 -172 1749 33
rect 4040 6 4069 58
rect 4121 6 4149 58
rect 4040 0 4149 6
rect 10358 189 10437 195
rect 10358 137 10371 189
rect 10423 137 10437 189
rect 10358 124 10437 137
rect 10358 72 10371 124
rect 10423 72 10437 124
rect 10358 58 10437 72
rect 10358 6 10371 58
rect 10423 6 10437 58
rect 10358 0 10437 6
rect 10790 -220 10831 195
<< via1 >>
rect 4227 3314 4279 3320
rect 4227 3280 4236 3314
rect 4236 3280 4270 3314
rect 4270 3280 4279 3314
rect 4227 3268 4279 3280
rect 4227 3242 4279 3254
rect 4227 3208 4236 3242
rect 4236 3208 4270 3242
rect 4270 3208 4279 3242
rect 4227 3202 4279 3208
rect 4327 3314 4379 3320
rect 4327 3280 4336 3314
rect 4336 3280 4370 3314
rect 4370 3280 4379 3314
rect 4327 3268 4379 3280
rect 4327 3242 4379 3254
rect 4327 3208 4336 3242
rect 4336 3208 4370 3242
rect 4370 3208 4379 3242
rect 4327 3202 4379 3208
rect 4483 3314 4535 3320
rect 4483 3280 4492 3314
rect 4492 3280 4526 3314
rect 4526 3280 4535 3314
rect 4483 3268 4535 3280
rect 4483 3242 4535 3254
rect 4483 3208 4492 3242
rect 4492 3208 4526 3242
rect 4526 3208 4535 3242
rect 4483 3202 4535 3208
rect 4585 3314 4637 3320
rect 4585 3280 4594 3314
rect 4594 3280 4628 3314
rect 4628 3280 4637 3314
rect 4585 3268 4637 3280
rect 4585 3242 4637 3254
rect 4585 3208 4594 3242
rect 4594 3208 4628 3242
rect 4628 3208 4637 3242
rect 4585 3202 4637 3208
rect 10069 3165 10121 3217
rect 4106 3054 4158 3106
rect 10069 3101 10121 3153
rect 10149 3167 10201 3219
rect 10149 3101 10201 3153
rect 10467 3167 10519 3219
rect 10467 3101 10519 3153
rect 10547 3165 10599 3217
rect 10547 3101 10599 3153
rect 4106 2979 4158 3031
rect 4106 2903 4158 2955
rect 10371 3001 10423 3053
rect 10371 2935 10423 2987
rect 10371 2869 10423 2921
rect 10208 2731 10260 2783
rect 10272 2731 10324 2783
rect 10467 2777 10519 2829
rect 12109 2783 12161 2835
rect 12173 2783 12225 2835
rect 10467 2713 10519 2765
rect 4333 2625 4385 2677
rect 4397 2625 4449 2677
rect 4489 2545 4541 2597
rect 4553 2545 4605 2597
rect 4233 2465 4285 2517
rect 4297 2465 4349 2517
rect 8334 2449 8386 2501
rect 8334 2385 8386 2437
rect 10278 2271 10330 2323
rect 10278 2207 10330 2259
rect 11402 2271 11454 2323
rect 11402 2207 11454 2259
rect 10003 1974 10055 2026
rect 10003 1910 10055 1962
rect 8334 1823 8386 1875
rect 8334 1759 8386 1811
rect 10371 1763 10423 1815
rect 6692 1673 6744 1725
rect 6756 1673 6808 1725
rect 10371 1688 10423 1740
rect 10371 1650 10423 1664
rect 9471 1593 9523 1645
rect 9535 1593 9587 1645
rect 10371 1616 10389 1650
rect 10389 1616 10423 1650
rect 10371 1612 10423 1616
rect 9933 1511 9985 1563
rect 9997 1511 10049 1563
rect 10192 1513 10244 1565
rect 10256 1513 10308 1565
rect 4726 1439 4778 1491
rect 4726 1375 4778 1427
rect 5712 1365 5764 1417
rect 5776 1365 5828 1417
rect 9547 1270 9599 1322
rect 9611 1270 9663 1322
rect 11102 1270 11154 1322
rect 11166 1270 11218 1322
rect 4069 137 4121 189
rect 4069 72 4121 124
rect 4069 6 4121 58
rect 10371 137 10423 189
rect 10371 72 10423 124
rect 10371 6 10423 58
<< metal2 >>
rect 4227 3320 4279 3326
rect 4227 3254 4279 3268
rect 4078 3106 4186 3112
rect 4078 3054 4106 3106
rect 4158 3054 4186 3106
rect 4078 3031 4186 3054
rect 4078 2979 4106 3031
rect 4158 2979 4186 3031
rect 4078 2955 4186 2979
rect 4078 2903 4106 2955
rect 4158 2903 4186 2955
tri 4040 2069 4078 2107 se
rect 4078 2069 4186 2903
rect 4227 2545 4279 3202
rect 4327 3320 4379 3326
rect 4327 3254 4379 3268
rect 4327 2677 4379 3202
rect 4483 3320 4535 3326
rect 4483 3254 4535 3268
tri 4379 2677 4413 2711 sw
rect 4327 2625 4333 2677
rect 4385 2625 4397 2677
rect 4449 2625 4455 2677
rect 4483 2625 4535 3202
rect 4585 3320 4695 3326
rect 4637 3268 4695 3320
rect 4585 3254 4695 3268
rect 4637 3202 4695 3254
rect 4585 3196 4695 3202
tri 4609 3165 4640 3196 ne
rect 4640 3165 4695 3196
tri 4640 3162 4643 3165 ne
rect 4643 2791 4695 3165
rect 10040 3217 10121 3223
rect 10040 3165 10069 3217
rect 10040 3153 10121 3165
rect 10040 3101 10069 3153
rect 10040 3095 10121 3101
tri 4695 2791 4704 2800 sw
rect 4643 2783 4704 2791
tri 4704 2783 4712 2791 sw
rect 4643 2778 4712 2783
tri 4643 2731 4690 2778 ne
rect 4690 2777 4712 2778
tri 4712 2777 4718 2783 sw
rect 4690 2731 4718 2777
tri 4718 2731 4764 2777 sw
rect 10040 2743 10092 3095
tri 10092 3066 10121 3095 nw
rect 10149 3219 10201 3245
rect 10547 3230 10916 3282
rect 10547 3225 10628 3230
tri 10628 3225 10633 3230 nw
tri 10830 3225 10835 3230 ne
rect 10835 3225 10916 3230
rect 10149 3153 10201 3167
rect 10149 2943 10201 3101
rect 10467 3219 10519 3225
rect 10467 3153 10519 3167
rect 10358 3053 10437 3059
rect 10358 3001 10371 3053
rect 10423 3001 10437 3053
rect 10358 2987 10437 3001
tri 10201 2943 10223 2965 sw
tri 10149 2935 10157 2943 ne
rect 10157 2935 10223 2943
tri 10223 2935 10231 2943 sw
rect 10358 2935 10371 2987
rect 10423 2935 10437 2987
tri 10157 2921 10171 2935 ne
rect 10171 2923 10231 2935
tri 10231 2923 10243 2935 sw
rect 10171 2921 10243 2923
tri 10171 2901 10191 2921 ne
rect 10191 2783 10243 2921
rect 10358 2921 10437 2935
rect 10358 2869 10371 2921
rect 10423 2869 10437 2921
tri 10243 2783 10277 2817 sw
tri 10040 2731 10052 2743 ne
rect 10052 2731 10092 2743
tri 10092 2731 10126 2765 sw
rect 10191 2731 10208 2783
rect 10260 2731 10272 2783
rect 10324 2731 10330 2783
tri 4690 2717 4704 2731 ne
rect 4704 2717 4764 2731
tri 4764 2717 4778 2731 sw
tri 4704 2713 4708 2717 ne
rect 4708 2713 4778 2717
tri 10052 2713 10070 2731 ne
rect 10070 2713 10126 2731
tri 10126 2713 10144 2731 sw
tri 10244 2713 10262 2731 ne
rect 10262 2713 10330 2731
tri 4708 2695 4726 2713 ne
tri 4535 2625 4541 2631 sw
rect 4483 2597 4541 2625
tri 4541 2597 4569 2625 sw
tri 4279 2545 4285 2551 sw
rect 4483 2545 4489 2597
rect 4541 2545 4553 2597
rect 4605 2545 4611 2597
rect 4227 2517 4285 2545
tri 4285 2517 4313 2545 sw
rect 4227 2465 4233 2517
rect 4285 2465 4297 2517
rect 4349 2465 4355 2517
rect 4040 2061 4186 2069
rect 4040 2026 4151 2061
tri 4151 2026 4186 2061 nw
rect 4040 189 4149 2026
tri 4149 2024 4151 2026 nw
rect 4726 1491 4778 2713
tri 10070 2693 10090 2713 ne
rect 10090 2693 10144 2713
tri 10144 2693 10164 2713 sw
tri 10262 2697 10278 2713 ne
tri 10090 2691 10092 2693 ne
rect 10092 2691 10164 2693
tri 10092 2635 10148 2691 ne
rect 10148 2635 10164 2691
rect 5285 2458 5357 2635
tri 10148 2619 10164 2635 ne
tri 10164 2619 10238 2693 sw
tri 10164 2597 10186 2619 ne
rect 8334 2501 8386 2507
rect 8334 2437 8386 2449
rect 6474 2136 6680 2188
tri 6658 2130 6664 2136 ne
rect 6664 2130 6680 2136
tri 6680 2130 6738 2188 sw
tri 6664 2114 6680 2130 ne
rect 6680 2114 6738 2130
tri 6680 2108 6686 2114 ne
rect 6686 1753 6738 2114
rect 8334 1875 8386 2385
rect 8334 1811 8386 1823
tri 6738 1753 6744 1759 sw
rect 8334 1753 8386 1759
rect 10003 2026 10055 2032
rect 10003 1962 10055 1974
rect 6686 1740 6744 1753
tri 6744 1740 6757 1753 sw
rect 6686 1725 6757 1740
tri 6757 1725 6772 1740 sw
rect 6686 1673 6692 1725
rect 6744 1673 6756 1725
rect 6808 1673 6814 1725
rect 9425 1593 9471 1645
rect 9523 1593 9535 1645
rect 9587 1593 9593 1645
tri 9507 1565 9535 1593 ne
rect 9535 1565 9593 1593
tri 9971 1565 10003 1597 se
rect 10003 1565 10055 1910
tri 9535 1563 9537 1565 ne
rect 9537 1563 9593 1565
tri 9969 1563 9971 1565 se
rect 9971 1563 10055 1565
tri 9537 1559 9541 1563 ne
rect 4726 1427 4778 1439
tri 5758 1417 5792 1451 sw
rect 4726 1369 4778 1375
rect 5706 1365 5712 1417
rect 5764 1365 5776 1417
rect 5828 1365 5834 1417
tri 5758 1331 5792 1365 nw
rect 9541 1322 9593 1563
rect 9927 1511 9933 1563
rect 9985 1511 9997 1563
rect 10049 1511 10055 1563
rect 10186 1565 10238 2619
rect 10278 2323 10330 2713
rect 10278 2259 10330 2271
rect 10278 2201 10330 2207
rect 10358 1815 10437 2869
rect 10467 2829 10519 3101
rect 10547 3223 10626 3225
tri 10626 3223 10628 3225 nw
tri 10835 3223 10837 3225 ne
rect 10837 3223 10916 3225
rect 10547 3217 10599 3223
tri 10599 3196 10626 3223 nw
tri 10837 3196 10864 3223 ne
rect 10864 3165 10916 3223
rect 10547 3153 10599 3165
rect 10547 3095 10599 3101
tri 12155 2835 12189 2869 sw
rect 12103 2783 12109 2835
rect 12161 2783 12173 2835
rect 12225 2783 12231 2835
rect 10467 2765 10519 2777
tri 12155 2749 12189 2783 nw
rect 10467 2707 10519 2713
rect 11402 2323 11454 2329
rect 11402 2259 11454 2271
rect 11402 2201 11454 2207
tri 11951 1836 11985 1870 sw
rect 10358 1763 10371 1815
rect 10423 1763 10437 1815
rect 10358 1740 10437 1763
rect 10358 1688 10371 1740
rect 10423 1688 10437 1740
tri 11917 1705 11951 1739 ne
rect 10358 1664 10437 1688
rect 10358 1612 10371 1664
rect 10423 1612 10437 1664
tri 10238 1565 10272 1599 sw
rect 10186 1513 10192 1565
rect 10244 1513 10256 1565
rect 10308 1513 10314 1565
tri 9593 1322 9627 1356 sw
rect 9541 1270 9547 1322
rect 9599 1270 9611 1322
rect 9663 1270 9669 1322
rect 10026 1208 10154 1241
rect 4040 137 4069 189
rect 4121 137 4149 189
rect 4040 124 4149 137
rect 4040 72 4069 124
rect 4121 72 4149 124
rect 4040 58 4149 72
rect 4040 6 4069 58
rect 4121 6 4149 58
rect 4040 0 4149 6
rect 10358 189 10437 1612
tri 11148 1322 11182 1356 sw
rect 11096 1270 11102 1322
rect 11154 1270 11166 1322
rect 11218 1270 11224 1322
tri 11148 1236 11182 1270 nw
rect 10358 137 10371 189
rect 10423 137 10437 189
rect 10358 124 10437 137
rect 10358 72 10371 124
rect 10423 72 10437 124
rect 10358 58 10437 72
rect 10358 6 10371 58
rect 10423 6 10437 58
rect 10358 0 10437 6
use sky130_fd_io__gpiov2_in_buf  sky130_fd_io__gpiov2_in_buf_0
timestamp 1683767628
transform 1 0 0 0 1 952
box -467 -1172 5758 3048
use sky130_fd_io__gpiov2_inbuf_lvinv_x1  sky130_fd_io__gpiov2_inbuf_lvinv_x1_0
timestamp 1683767628
transform -1 0 10609 0 1 2831
box 0 0 359 1066
use sky130_fd_io__gpiov2_inbuf_lvinv_x1  sky130_fd_io__gpiov2_inbuf_lvinv_x1_1
timestamp 1683767628
transform 1 0 10059 0 1 2831
box 0 0 359 1066
use sky130_fd_io__gpiov2_ipath_hvls  sky130_fd_io__gpiov2_ipath_hvls_0
timestamp 1683767628
transform -1 0 8860 0 1 -51
box 536 -169 4076 4051
use sky130_fd_io__gpiov2_ipath_lvls  sky130_fd_io__gpiov2_ipath_lvls_0
timestamp 1683767628
transform -1 0 12999 0 1 471
box 74 -691 2336 3529
use sky130_fd_io__gpiov2_vcchib_in_buf  sky130_fd_io__gpiov2_vcchib_in_buf_0
timestamp 1683767628
transform 1 0 8210 0 1 355
box 114 -575 2586 3645
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1683767628
transform 1 0 4344 0 1 2873
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_1
timestamp 1683767628
transform -1 0 4526 0 1 2873
box 107 226 240 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1683767628
transform -1 0 10706 0 1 1582
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_1
timestamp 1683767628
transform 1 0 10524 0 1 1582
box 107 226 460 873
<< labels >>
flabel metal1 s 265 1382 375 1423 3 FreeSans 200 0 0 0 VTRIP_SEL_H_N
port 2 nsew
flabel metal1 s 11495 3762 12100 3985 3 FreeSans 200 0 0 0 VCCHIB
port 3 nsew
flabel metal1 s 10519 1934 10604 1965 3 FreeSans 200 0 0 0 ENABLE_VDDIO_LV
port 4 nsew
flabel metal1 s 99 2628 266 2672 3 FreeSans 200 0 0 0 MODE_NORMAL_N
port 5 nsew
flabel metal1 s 1179 -172 1749 33 3 FreeSans 200 0 0 0 VSSD
port 6 nsew
flabel metal1 s 954 3782 1636 3954 3 FreeSans 200 0 0 0 VDDIO_Q
port 7 nsew
flabel metal1 s 12230 1946 12377 1995 3 FreeSans 200 0 0 0 IBUFMUX_OUT
port 8 nsew
flabel metal1 s 397 2393 483 2427 3 FreeSans 200 0 0 0 IN_VT
port 9 nsew
flabel metal1 s 384 1293 476 1325 3 FreeSans 200 0 0 0 IN_H
port 10 nsew
flabel metal1 s 265 2069 398 2104 3 FreeSans 200 0 0 0 VTRIP_SEL_H
port 11 nsew
flabel metal1 s 99 2552 241 2589 3 FreeSans 200 0 0 0 MODE_VCCHIB_N
port 12 nsew
flabel metal2 s 5285 2458 5357 2635 3 FreeSans 200 0 0 0 IBUFMUX_OUT_H
port 13 nsew
<< properties >>
string GDS_END 3703954
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3676042
<< end >>
