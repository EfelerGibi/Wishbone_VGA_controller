magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -66 377 834 897
<< pwell >>
rect -26 -43 794 43
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 831 768 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
rect 0 791 768 797
rect 0 689 768 763
rect 0 51 768 125
rect 0 17 768 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -23 768 -17
<< labels >>
rlabel metal1 s 0 51 768 125 6 VGND
port 1 nsew ground bidirectional
rlabel metal1 s 0 -23 768 23 8 VNB
port 2 nsew ground bidirectional
rlabel pwell s -26 -43 794 43 8 VNB
port 2 nsew ground bidirectional
rlabel metal1 s 0 791 768 837 6 VPB
port 3 nsew power bidirectional
rlabel nwell s -66 377 834 897 6 VPB
port 3 nsew power bidirectional
rlabel metal1 s 0 689 768 763 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 768 814
string LEFclass CORE SPACER
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 87736
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 82668
<< end >>
