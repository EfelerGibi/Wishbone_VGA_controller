magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 1 21 911 203
rect 29 -17 63 21
<< scnmos >>
rect 84 47 114 177
rect 170 47 200 177
rect 256 47 286 177
rect 342 47 372 177
rect 540 47 570 177
rect 626 47 656 177
rect 712 47 742 177
rect 798 47 828 177
<< scpmoshvt >>
rect 84 297 114 497
rect 170 297 200 497
rect 256 297 286 497
rect 342 297 372 497
rect 540 297 570 497
rect 626 297 656 497
rect 712 297 742 497
rect 798 297 828 497
<< ndiff >>
rect 27 89 84 177
rect 27 55 39 89
rect 73 55 84 89
rect 27 47 84 55
rect 114 169 170 177
rect 114 135 125 169
rect 159 135 170 169
rect 114 47 170 135
rect 200 158 256 177
rect 200 124 211 158
rect 245 124 256 158
rect 200 89 256 124
rect 200 55 211 89
rect 245 55 256 89
rect 200 47 256 55
rect 286 165 342 177
rect 286 131 297 165
rect 331 131 342 165
rect 286 47 342 131
rect 372 89 429 177
rect 372 55 383 89
rect 417 55 429 89
rect 372 47 429 55
rect 483 89 540 177
rect 483 55 495 89
rect 529 55 540 89
rect 483 47 540 55
rect 570 165 626 177
rect 570 131 581 165
rect 615 131 626 165
rect 570 47 626 131
rect 656 89 712 177
rect 656 55 667 89
rect 701 55 712 89
rect 656 47 712 55
rect 742 153 798 177
rect 742 119 753 153
rect 787 119 798 153
rect 742 47 798 119
rect 828 89 885 177
rect 828 55 839 89
rect 873 55 885 89
rect 828 47 885 55
<< pdiff >>
rect 31 485 84 497
rect 31 451 39 485
rect 73 451 84 485
rect 31 297 84 451
rect 114 477 170 497
rect 114 443 125 477
rect 159 443 170 477
rect 114 381 170 443
rect 114 347 125 381
rect 159 347 170 381
rect 114 297 170 347
rect 200 485 256 497
rect 200 451 211 485
rect 245 451 256 485
rect 200 417 256 451
rect 200 383 211 417
rect 245 383 256 417
rect 200 297 256 383
rect 286 477 342 497
rect 286 443 297 477
rect 331 443 342 477
rect 286 386 342 443
rect 286 352 297 386
rect 331 352 342 386
rect 286 297 342 352
rect 372 485 425 497
rect 372 451 383 485
rect 417 451 425 485
rect 372 417 425 451
rect 372 383 383 417
rect 417 383 425 417
rect 372 297 425 383
rect 487 477 540 497
rect 487 443 495 477
rect 529 443 540 477
rect 487 297 540 443
rect 570 425 626 497
rect 570 391 581 425
rect 615 391 626 425
rect 570 357 626 391
rect 570 323 581 357
rect 615 323 626 357
rect 570 297 626 323
rect 656 477 712 497
rect 656 443 667 477
rect 701 443 712 477
rect 656 382 712 443
rect 656 348 667 382
rect 701 348 712 382
rect 656 297 712 348
rect 742 485 798 497
rect 742 451 753 485
rect 787 451 798 485
rect 742 407 798 451
rect 742 373 753 407
rect 787 373 798 407
rect 742 297 798 373
rect 828 477 881 497
rect 828 443 839 477
rect 873 443 881 477
rect 828 409 881 443
rect 828 375 839 409
rect 873 375 881 409
rect 828 297 881 375
<< ndiffc >>
rect 39 55 73 89
rect 125 135 159 169
rect 211 124 245 158
rect 211 55 245 89
rect 297 131 331 165
rect 383 55 417 89
rect 495 55 529 89
rect 581 131 615 165
rect 667 55 701 89
rect 753 119 787 153
rect 839 55 873 89
<< pdiffc >>
rect 39 451 73 485
rect 125 443 159 477
rect 125 347 159 381
rect 211 451 245 485
rect 211 383 245 417
rect 297 443 331 477
rect 297 352 331 386
rect 383 451 417 485
rect 383 383 417 417
rect 495 443 529 477
rect 581 391 615 425
rect 581 323 615 357
rect 667 443 701 477
rect 667 348 701 382
rect 753 451 787 485
rect 753 373 787 407
rect 839 443 873 477
rect 839 375 873 409
<< poly >>
rect 84 497 114 523
rect 170 497 200 523
rect 256 497 286 523
rect 342 497 372 523
rect 540 497 570 523
rect 626 497 656 523
rect 712 497 742 523
rect 798 497 828 523
rect 84 265 114 297
rect 170 265 200 297
rect 256 265 286 297
rect 342 265 372 297
rect 540 265 570 297
rect 626 265 656 297
rect 712 265 742 297
rect 798 265 828 297
rect 21 249 200 265
rect 21 215 31 249
rect 65 215 200 249
rect 21 199 200 215
rect 242 249 372 265
rect 242 215 252 249
rect 286 215 320 249
rect 354 215 372 249
rect 242 199 372 215
rect 539 249 661 265
rect 539 215 549 249
rect 583 215 617 249
rect 651 215 661 249
rect 539 199 661 215
rect 707 249 829 265
rect 707 215 717 249
rect 751 215 785 249
rect 819 215 829 249
rect 707 199 829 215
rect 84 177 114 199
rect 170 177 200 199
rect 256 177 286 199
rect 342 177 372 199
rect 540 177 570 199
rect 626 177 656 199
rect 712 177 742 199
rect 798 177 828 199
rect 84 21 114 47
rect 170 21 200 47
rect 256 21 286 47
rect 342 21 372 47
rect 540 21 570 47
rect 626 21 656 47
rect 712 21 742 47
rect 798 21 828 47
<< polycont >>
rect 31 215 65 249
rect 252 215 286 249
rect 320 215 354 249
rect 549 215 583 249
rect 617 215 651 249
rect 717 215 751 249
rect 785 215 819 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 23 485 75 527
rect 23 451 39 485
rect 73 451 75 485
rect 23 435 75 451
rect 109 477 161 493
rect 109 443 125 477
rect 159 443 161 477
rect 17 249 75 394
rect 17 215 31 249
rect 65 215 75 249
rect 17 199 75 215
rect 109 381 161 443
rect 195 485 261 527
rect 195 451 211 485
rect 245 451 261 485
rect 195 417 261 451
rect 195 383 211 417
rect 245 383 261 417
rect 295 477 333 493
rect 295 443 297 477
rect 331 443 333 477
rect 295 386 333 443
rect 109 347 125 381
rect 159 347 161 381
rect 109 342 161 347
rect 295 352 297 386
rect 331 352 333 386
rect 367 485 433 527
rect 367 451 383 485
rect 417 451 433 485
rect 367 417 433 451
rect 479 477 703 493
rect 479 443 495 477
rect 529 459 667 477
rect 529 443 531 459
rect 479 420 531 443
rect 665 443 667 459
rect 701 443 703 477
rect 367 383 383 417
rect 417 383 433 417
rect 565 391 581 425
rect 615 391 631 425
rect 295 342 333 352
rect 565 357 631 391
rect 565 342 581 357
rect 109 323 581 342
rect 615 323 631 357
rect 109 308 631 323
rect 665 382 703 443
rect 665 348 667 382
rect 701 348 703 382
rect 737 485 803 527
rect 737 451 753 485
rect 787 451 803 485
rect 737 407 803 451
rect 737 373 753 407
rect 787 373 803 407
rect 837 477 889 493
rect 837 443 839 477
rect 873 443 889 477
rect 837 409 889 443
rect 837 375 839 409
rect 873 375 889 409
rect 665 339 703 348
rect 837 339 889 375
rect 109 169 175 308
rect 665 305 889 339
rect 209 249 381 273
rect 209 215 252 249
rect 286 215 320 249
rect 354 215 381 249
rect 473 249 667 271
rect 712 249 891 259
rect 473 215 549 249
rect 583 215 617 249
rect 651 215 667 249
rect 701 215 717 249
rect 751 215 785 249
rect 819 215 891 249
rect 109 135 125 169
rect 159 135 175 169
rect 109 134 175 135
rect 209 158 247 178
rect 209 124 211 158
rect 245 124 247 158
rect 281 165 789 169
rect 281 131 297 165
rect 331 131 581 165
rect 615 153 789 165
rect 823 153 891 215
rect 615 131 753 153
rect 281 127 753 131
rect 209 93 247 124
rect 751 119 753 127
rect 787 119 789 153
rect 751 103 789 119
rect 209 89 433 93
rect 19 55 39 89
rect 73 55 211 89
rect 245 55 383 89
rect 417 55 433 89
rect 19 51 433 55
rect 479 55 495 89
rect 529 55 545 89
rect 479 17 545 55
rect 651 55 667 89
rect 701 55 717 89
rect 651 17 717 55
rect 823 55 839 89
rect 873 55 889 89
rect 823 17 889 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel locali s 857 153 891 187 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 121 153 155 187 0 FreeSans 400 0 0 0 Y
port 9 nsew signal output
flabel locali s 29 289 63 323 0 FreeSans 400 0 0 0 C1
port 4 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o211ai_2
rlabel metal1 s 0 -48 920 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 920 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 783804
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 776408
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 4.600 0.000 
<< end >>
