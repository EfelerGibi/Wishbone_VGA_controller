magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< metal2 >>
rect 9499 -407 14279 -259
rect 14579 -407 14979 -211
rect 19478 -407 24258 -259
<< metal3 >>
tri 0 27305 6919 34224 se
rect 6919 27305 9579 34224
rect 0 22525 9579 27305
rect 0 2730 4307 22525
tri 4307 22327 4505 22525 nw
tri 4897 22327 5095 22525 ne
rect 5095 22327 9579 22525
tri 5095 22325 5097 22327 ne
rect 5097 21630 9579 22327
rect 5096 16548 9579 21630
tri 5093 2927 5096 2930 se
rect 5096 2927 8904 16548
tri 8904 16348 9104 16548 nw
tri 9299 16348 9499 16548 ne
rect 9499 16348 9579 16548
rect 24146 27295 26838 34257
tri 26838 27295 33800 34257 sw
rect 24146 22525 33800 27295
rect 24146 21725 28705 22525
tri 28705 22325 28905 22525 nw
tri 29296 22325 29496 22525 ne
rect 24146 16548 28704 21725
rect 24146 16348 24258 16548
tri 24258 16348 24458 16548 nw
tri 24696 16348 24896 16548 ne
tri 4307 2730 4504 2927 sw
tri 4896 2730 5093 2927 se
rect 5093 2730 8904 2927
tri 8904 2730 9104 2930 sw
tri 9299 2730 9499 2930 se
rect 9499 2730 9579 2930
rect 0 -16 9579 2730
rect 24146 2730 24258 2930
tri 24258 2730 24458 2930 sw
tri 24696 2730 24896 2930 se
rect 24896 2730 28704 16548
tri 28704 2730 28904 2930 sw
tri 29296 2730 29496 2930 se
rect 29496 2730 33800 22525
rect 24146 -16 33800 2730
rect 0 -407 14279 -16
rect 14579 -407 16779 -259
rect 16978 -407 19178 -89
rect 19478 -407 33800 -16
<< metal4 >>
rect 0 34750 254 39593
rect 33546 34750 33800 39593
rect 0 13600 254 18593
rect 33546 13600 33800 18593
rect 0 12410 254 13300
rect 33546 12410 33800 13300
rect 0 11240 254 12130
rect 33546 11240 33800 12130
rect 0 10874 254 10940
rect 33546 10874 33800 10940
rect 0 10218 254 10814
rect 33546 10218 33800 10814
rect 0 9922 254 10158
rect 33546 9922 33800 10158
rect 0 9266 254 9862
rect 33546 9266 33800 9862
rect 0 9140 254 9206
rect 33546 9140 33800 9206
rect 0 7910 254 8840
rect 33546 7910 33800 8840
rect 0 6940 254 7630
rect 33546 6940 33800 7630
rect 0 5970 254 6660
rect 33546 5970 33800 6660
rect 0 4760 254 5690
rect 33546 4760 33800 5690
rect 0 3550 254 4480
rect 33546 3550 33800 4480
rect 0 2580 254 3270
rect 33546 2580 33800 3270
rect 0 1370 254 2300
rect 33546 1370 33800 2300
rect 0 0 254 1090
rect 33546 0 33800 1090
<< metal5 >>
rect 0 34750 254 39593
rect 33546 34750 33800 39593
rect 16729 27458 16994 28780
rect 0 13600 254 18590
rect 33546 13600 33800 18590
rect 0 12430 254 13280
rect 33546 12430 33800 13280
rect 0 11260 254 12110
rect 33546 11260 33800 12110
rect 0 9140 254 10940
rect 33546 9140 33800 10940
rect 0 7930 254 8820
rect 33546 7930 33800 8820
rect 0 6960 254 7610
rect 33546 6960 33800 7610
rect 0 5990 254 6640
rect 33546 5990 33800 6640
rect 0 4780 254 5670
rect 33546 4780 33800 5670
rect 0 3570 254 4460
rect 33546 3570 33800 4460
rect 0 2600 254 3250
rect 33546 2600 33800 3250
rect 0 1390 254 2280
rect 33546 1390 33800 2280
rect 0 20 254 1070
rect 33546 20 33800 1070
use sky130_ef_io__com_bus_slice_1um  sky130_ef_io__com_bus_slice_1um_0
timestamp 1683767628
transform 1 0 33400 0 1 0
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  sky130_ef_io__com_bus_slice_1um_1
timestamp 1683767628
transform 1 0 33600 0 1 0
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  sky130_ef_io__com_bus_slice_1um_2
timestamp 1683767628
transform 1 0 0 0 1 0
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  sky130_ef_io__com_bus_slice_1um_3
timestamp 1683767628
transform 1 0 200 0 1 0
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_0
timestamp 1683767628
transform 1 0 32400 0 1 0
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_1
timestamp 1683767628
transform 1 0 400 0 1 0
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_0
timestamp 1683767628
transform 1 0 24400 0 1 0
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_1
timestamp 1683767628
transform 1 0 28400 0 1 0
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_2
timestamp 1683767628
transform 1 0 1400 0 1 0
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_3
timestamp 1683767628
transform 1 0 5400 0 1 0
box 0 0 4000 39593
use sky130_fd_io__top_power_hvc_wpadv2  sky130_fd_io__top_power_hvc_wpadv2_1
timestamp 1683767628
transform 1 0 9400 0 1 -407
box 0 0 15000 40000
<< labels >>
flabel metal4 s 0 10218 254 10814 3 FreeSans 650 0 0 0 AMUXBUS_A
port 1 nsew
flabel metal4 s 33546 10218 33800 10814 3 FreeSans 650 180 0 0 AMUXBUS_A
port 1 nsew
flabel metal4 s 0 9266 254 9862 3 FreeSans 650 0 0 0 AMUXBUS_B
port 2 nsew
flabel metal4 s 33546 9266 33800 9862 3 FreeSans 650 180 0 0 AMUXBUS_B
port 2 nsew
flabel metal3 s 16978 -407 19178 -89 0 FreeSans 2500 0 0 0 DRN_HVC
port 3 nsew
flabel metal2 s 19478 -407 24258 -259 2 FreeSans 2500 90 0 0 DRN_HVC
port 3 nsew
flabel metal3 s 19478 -407 33757 -16 0 FreeSans 2500 0 0 0 P_CORE
port 4 nsew
flabel metal3 s 0 -407 14279 -16 0 FreeSans 2500 0 0 0 P_CORE
port 4 nsew
flabel metal5 s 16729 27458 16994 28780 0 FreeSans 2500 0 0 0 P_PAD
port 5 nsew
flabel metal3 s 14579 -407 16779 -259 2 FreeSans 2500 90 0 0 SRC_BDY_HVC
port 6 nsew
flabel metal2 s 9499 -407 14279 -259 2 FreeSans 2500 90 0 0 SRC_BDY_HVC
port 6 nsew
flabel metal4 s 0 6940 254 7630 3 FreeSans 650 0 0 0 VSSA
port 8 nsew
flabel metal4 s 0 10874 254 10940 3 FreeSans 650 0 0 0 VSSA
port 8 nsew
flabel metal4 s 0 9922 254 10158 3 FreeSans 650 0 0 0 VSSA
port 8 nsew
flabel metal4 s 0 9140 254 9206 3 FreeSans 650 0 0 0 VSSA
port 8 nsew
flabel metal5 s 0 6961 254 7610 3 FreeSans 650 0 0 0 VSSA
port 8 nsew
flabel metal5 s 0 9140 254 10940 3 FreeSans 650 0 0 0 VSSA
port 8 nsew
flabel metal4 s 33546 6940 33800 7630 3 FreeSans 650 180 0 0 VSSA
port 8 nsew
flabel metal4 s 33546 9140 33800 9206 3 FreeSans 650 180 0 0 VSSA
port 8 nsew
flabel metal4 s 33546 10874 33800 10940 3 FreeSans 650 180 0 0 VSSA
port 8 nsew
flabel metal4 s 33546 9922 33800 10158 3 FreeSans 650 180 0 0 VSSA
port 8 nsew
flabel metal5 s 33546 6961 33800 7610 3 FreeSans 650 180 0 0 VSSA
port 8 nsew
flabel metal5 s 33546 9140 33800 10940 3 FreeSans 650 180 0 0 VSSA
port 8 nsew
flabel metal4 s 0 2580 193 3270 3 FreeSans 650 0 0 0 VDDA
port 9 nsew
flabel metal5 s 0 2600 193 3250 3 FreeSans 650 0 0 0 VDDA
port 9 nsew
flabel metal4 s 33607 2580 33800 3270 3 FreeSans 650 180 0 0 VDDA
port 9 nsew
flabel metal5 s 33607 2600 33800 3250 3 FreeSans 650 180 0 0 VDDA
port 9 nsew
flabel metal4 s 0 5970 254 6660 3 FreeSans 650 0 0 0 VSWITCH
port 10 nsew
flabel metal5 s 0 5990 254 6640 3 FreeSans 650 0 0 0 VSWITCH
port 10 nsew
flabel metal4 s 33546 5970 33800 6660 3 FreeSans 650 180 0 0 VSWITCH
port 10 nsew
flabel metal5 s 33546 5990 33800 6640 3 FreeSans 650 180 0 0 VSWITCH
port 10 nsew
flabel metal4 s 0 12410 254 13300 3 FreeSans 650 0 0 0 VDDIO_Q
port 11 nsew
flabel metal5 s 0 12430 254 13280 3 FreeSans 650 0 0 0 VDDIO_Q
port 11 nsew
flabel metal4 s 33546 12410 33800 13300 3 FreeSans 650 180 0 0 VDDIO_Q
port 11 nsew
flabel metal5 s 33546 12430 33800 13280 3 FreeSans 650 180 0 0 VDDIO_Q
port 11 nsew
flabel metal4 s 0 0 254 1090 3 FreeSans 650 0 0 0 VCCHIB
port 12 nsew
flabel metal5 s 0 20 254 1070 3 FreeSans 650 0 0 0 VCCHIB
port 12 nsew
flabel metal4 s 33546 0 33800 1090 3 FreeSans 650 180 0 0 VCCHIB
port 12 nsew
flabel metal5 s 33546 20 33800 1070 3 FreeSans 650 180 0 0 VCCHIB
port 12 nsew
flabel metal4 s 0 13600 254 18593 3 FreeSans 650 0 0 0 VDDIO
port 13 nsew
flabel metal4 s 0 3550 254 4480 3 FreeSans 650 0 0 0 VDDIO
port 13 nsew
flabel metal5 s 0 3570 254 4460 3 FreeSans 650 0 0 0 VDDIO
port 13 nsew
flabel metal5 s 0 13600 254 18590 3 FreeSans 650 0 0 0 VDDIO
port 13 nsew
flabel metal4 s 33546 13600 33800 18593 3 FreeSans 650 180 0 0 VDDIO
port 13 nsew
flabel metal4 s 33546 3550 33800 4480 3 FreeSans 650 180 0 0 VDDIO
port 13 nsew
flabel metal5 s 33546 3570 33800 4460 3 FreeSans 650 180 0 0 VDDIO
port 13 nsew
flabel metal5 s 33546 13600 33800 18590 3 FreeSans 650 180 0 0 VDDIO
port 13 nsew
flabel metal4 s 0 1370 254 2300 3 FreeSans 650 0 0 0 VCCD
port 14 nsew
flabel metal5 s 0 1390 254 2280 3 FreeSans 650 0 0 0 VCCD
port 14 nsew
flabel metal4 s 33546 1370 33800 2300 3 FreeSans 650 180 0 0 VCCD
port 14 nsew
flabel metal5 s 33546 1390 33800 2280 3 FreeSans 650 180 0 0 VCCD
port 14 nsew
flabel metal4 s 0 4760 254 5690 3 FreeSans 650 0 0 0 VSSIO
port 15 nsew
flabel metal4 s 0 34750 254 39593 3 FreeSans 650 0 0 0 VSSIO
port 15 nsew
flabel metal5 s 0 4780 254 5670 3 FreeSans 650 0 0 0 VSSIO
port 15 nsew
flabel metal4 s 127 37914 127 37914 3 FreeSans 650 0 0 0 VSSIO
flabel metal4 s 127 37925 127 37925 3 FreeSans 650 0 0 0 VSSIO
flabel metal4 s 33546 34750 33800 39593 3 FreeSans 650 180 0 0 VSSIO
port 15 nsew
flabel metal4 s 33546 4760 33800 5690 3 FreeSans 650 180 0 0 VSSIO
port 15 nsew
flabel metal5 s 33546 4780 33800 5670 3 FreeSans 650 180 0 0 VSSIO
port 15 nsew
flabel metal4 s 33673 37914 33673 37914 3 FreeSans 650 180 0 0 VSSIO
flabel metal4 s 33673 37925 33673 37925 3 FreeSans 650 180 0 0 VSSIO
flabel metal4 s 0 7910 254 8840 3 FreeSans 650 0 0 0 VSSD
port 16 nsew
flabel metal5 s 0 7930 254 8820 3 FreeSans 650 0 0 0 VSSD
port 16 nsew
flabel metal4 s 33546 7910 33800 8840 3 FreeSans 650 180 0 0 VSSD
port 16 nsew
flabel metal5 s 33546 7930 33800 8820 3 FreeSans 650 180 0 0 VSSD
port 16 nsew
flabel metal4 s 0 11240 254 12130 3 FreeSans 650 0 0 0 VSSIO_Q
port 17 nsew
flabel metal5 s 0 11260 254 12110 3 FreeSans 650 0 0 0 VSSIO_Q
port 17 nsew
flabel metal4 s 33546 11240 33800 12130 3 FreeSans 650 180 0 0 VSSIO_Q
port 17 nsew
flabel metal5 s 33546 11260 33800 12110 3 FreeSans 650 180 0 0 VSSIO_Q
port 17 nsew
<< properties >>
string FIXED_BBOX 0 0 33800 39593
string GDS_END 3673392
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_START 3656272
<< end >>
