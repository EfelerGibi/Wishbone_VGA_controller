* NGSPICE file created from sky130_fd_pr__rf_pnp_05v5_W3p40L3p40.ext - technology: sky130B

.subckt sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 Emitter Collector Base
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0
**devattr s=37813,302
.ends

