magic
tech sky130B
timestamp 1683767628
<< properties >>
string GDS_END 12231328
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 12231004
<< end >>
