magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -36 679 8292 1471
<< locali >>
rect 0 1397 8256 1431
rect 64 636 98 702
rect 196 652 449 686
rect 547 653 817 687
rect 919 674 1293 708
rect 1609 690 2093 724
rect 2858 690 3757 724
rect 5911 690 5945 724
rect 919 670 953 674
rect 0 -17 8256 17
use sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6  sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_0
timestamp 1683767628
transform 1 0 368 0 1 0
box -36 -17 404 1471
use sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6  sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_1
timestamp 1683767628
transform 1 0 0 0 1 0
box -36 -17 404 1471
use sky130_sram_1kbyte_1rw1r_32x256_8_pinv_7  sky130_sram_1kbyte_1rw1r_32x256_8_pinv_7_0
timestamp 1683767628
transform 1 0 736 0 1 0
box -36 -17 512 1471
use sky130_sram_1kbyte_1rw1r_32x256_8_pinv_8  sky130_sram_1kbyte_1rw1r_32x256_8_pinv_8_0
timestamp 1683767628
transform 1 0 1212 0 1 0
box -36 -17 836 1471
use sky130_sram_1kbyte_1rw1r_32x256_8_pinv_9  sky130_sram_1kbyte_1rw1r_32x256_8_pinv_9_0
timestamp 1683767628
transform 1 0 2012 0 1 0
box -36 -17 1700 1471
use sky130_sram_1kbyte_1rw1r_32x256_8_pinv_10  sky130_sram_1kbyte_1rw1r_32x256_8_pinv_10_0
timestamp 1683767628
transform 1 0 3676 0 1 0
box -36 -17 4616 1471
<< labels >>
rlabel locali s 5928 707 5928 707 4 Z
rlabel locali s 81 669 81 669 4 A
rlabel locali s 4128 0 4128 0 4 gnd
rlabel locali s 4128 1414 4128 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 8256 1414
string GDS_END 6275200
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 6273314
<< end >>
