magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 1 21 1287 203
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 527 47 557 177
rect 599 47 629 177
rect 718 47 748 177
rect 804 47 834 177
rect 898 47 928 177
rect 1006 47 1036 177
rect 1092 47 1122 177
rect 1178 47 1208 177
<< scpmoshvt >>
rect 157 297 187 497
rect 243 297 273 497
rect 329 297 359 497
rect 415 297 445 497
rect 501 297 531 497
rect 632 297 662 497
rect 718 297 748 497
rect 826 297 856 497
rect 920 297 950 497
rect 1006 297 1036 497
rect 1092 297 1122 497
rect 1178 297 1208 497
<< ndiff >>
rect 27 93 79 177
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 101 163 177
rect 109 67 119 101
rect 153 67 163 101
rect 109 47 163 67
rect 193 89 247 177
rect 193 55 203 89
rect 237 55 247 89
rect 193 47 247 55
rect 277 101 331 177
rect 277 67 287 101
rect 321 67 331 101
rect 277 47 331 67
rect 361 93 420 177
rect 361 59 371 93
rect 405 59 420 93
rect 361 47 420 59
rect 474 93 527 177
rect 474 59 482 93
rect 516 59 527 93
rect 474 47 527 59
rect 557 47 599 177
rect 629 163 718 177
rect 629 129 654 163
rect 688 129 718 163
rect 629 47 718 129
rect 748 47 804 177
rect 834 169 898 177
rect 834 135 850 169
rect 884 135 898 169
rect 834 101 898 135
rect 834 67 850 101
rect 884 67 898 101
rect 834 47 898 67
rect 928 89 1006 177
rect 928 55 947 89
rect 981 55 1006 89
rect 928 47 1006 55
rect 1036 157 1092 177
rect 1036 123 1047 157
rect 1081 123 1092 157
rect 1036 89 1092 123
rect 1036 55 1047 89
rect 1081 55 1092 89
rect 1036 47 1092 55
rect 1122 89 1178 177
rect 1122 55 1133 89
rect 1167 55 1178 89
rect 1122 47 1178 55
rect 1208 161 1261 177
rect 1208 127 1219 161
rect 1253 127 1261 161
rect 1208 93 1261 127
rect 1208 59 1219 93
rect 1253 59 1261 93
rect 1208 47 1261 59
<< pdiff >>
rect 104 485 157 497
rect 104 451 112 485
rect 146 451 157 485
rect 104 408 157 451
rect 104 374 112 408
rect 146 374 157 408
rect 104 297 157 374
rect 187 477 243 497
rect 187 443 198 477
rect 232 443 243 477
rect 187 386 243 443
rect 187 352 198 386
rect 232 352 243 386
rect 187 297 243 352
rect 273 485 329 497
rect 273 451 284 485
rect 318 451 329 485
rect 273 408 329 451
rect 273 374 284 408
rect 318 374 329 408
rect 273 297 329 374
rect 359 477 415 497
rect 359 443 370 477
rect 404 443 415 477
rect 359 386 415 443
rect 359 352 370 386
rect 404 352 415 386
rect 359 297 415 352
rect 445 481 501 497
rect 445 447 456 481
rect 490 447 501 481
rect 445 297 501 447
rect 531 477 632 497
rect 531 443 562 477
rect 596 443 632 477
rect 531 297 632 443
rect 662 489 718 497
rect 662 455 673 489
rect 707 455 718 489
rect 662 297 718 455
rect 748 477 826 497
rect 748 443 773 477
rect 807 443 826 477
rect 748 297 826 443
rect 856 489 920 497
rect 856 455 867 489
rect 901 455 920 489
rect 856 297 920 455
rect 950 297 1006 497
rect 1036 489 1092 497
rect 1036 455 1047 489
rect 1081 455 1092 489
rect 1036 421 1092 455
rect 1036 387 1047 421
rect 1081 387 1092 421
rect 1036 297 1092 387
rect 1122 297 1178 497
rect 1208 485 1261 497
rect 1208 451 1219 485
rect 1253 451 1261 485
rect 1208 417 1261 451
rect 1208 383 1219 417
rect 1253 383 1261 417
rect 1208 297 1261 383
<< ndiffc >>
rect 35 59 69 93
rect 119 67 153 101
rect 203 55 237 89
rect 287 67 321 101
rect 371 59 405 93
rect 482 59 516 93
rect 654 129 688 163
rect 850 135 884 169
rect 850 67 884 101
rect 947 55 981 89
rect 1047 123 1081 157
rect 1047 55 1081 89
rect 1133 55 1167 89
rect 1219 127 1253 161
rect 1219 59 1253 93
<< pdiffc >>
rect 112 451 146 485
rect 112 374 146 408
rect 198 443 232 477
rect 198 352 232 386
rect 284 451 318 485
rect 284 374 318 408
rect 370 443 404 477
rect 370 352 404 386
rect 456 447 490 481
rect 562 443 596 477
rect 673 455 707 489
rect 773 443 807 477
rect 867 455 901 489
rect 1047 455 1081 489
rect 1047 387 1081 421
rect 1219 451 1253 485
rect 1219 383 1253 417
<< poly >>
rect 157 497 187 523
rect 243 497 273 523
rect 329 497 359 523
rect 415 497 445 523
rect 501 497 531 523
rect 632 497 662 523
rect 718 497 748 523
rect 826 497 856 523
rect 920 497 950 523
rect 1006 497 1036 523
rect 1092 497 1122 523
rect 1178 497 1208 523
rect 157 265 187 297
rect 243 265 273 297
rect 329 265 359 297
rect 415 265 445 297
rect 501 265 531 297
rect 632 265 662 297
rect 718 265 748 297
rect 826 265 856 297
rect 920 265 950 297
rect 1006 265 1036 297
rect 1092 265 1122 297
rect 1178 265 1208 297
rect 79 249 445 265
rect 79 215 123 249
rect 157 215 191 249
rect 225 215 259 249
rect 293 215 327 249
rect 361 215 395 249
rect 429 215 445 249
rect 79 199 445 215
rect 498 249 557 265
rect 498 215 508 249
rect 542 215 557 249
rect 498 199 557 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 331 177 361 199
rect 527 177 557 199
rect 599 249 748 265
rect 599 215 630 249
rect 664 215 698 249
rect 732 215 748 249
rect 599 199 748 215
rect 790 249 856 265
rect 790 215 806 249
rect 840 215 856 249
rect 790 199 856 215
rect 898 249 964 265
rect 898 215 914 249
rect 948 215 964 249
rect 898 199 964 215
rect 1006 249 1136 265
rect 1006 215 1022 249
rect 1056 215 1090 249
rect 1124 215 1136 249
rect 1006 199 1136 215
rect 1178 249 1258 265
rect 1178 215 1200 249
rect 1234 215 1258 249
rect 1178 199 1258 215
rect 599 177 629 199
rect 718 177 748 199
rect 804 177 834 199
rect 898 177 928 199
rect 1006 177 1036 199
rect 1092 177 1122 199
rect 1178 177 1208 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 527 21 557 47
rect 599 21 629 47
rect 718 21 748 47
rect 804 21 834 47
rect 898 21 928 47
rect 1006 21 1036 47
rect 1092 21 1122 47
rect 1178 21 1208 47
<< polycont >>
rect 123 215 157 249
rect 191 215 225 249
rect 259 215 293 249
rect 327 215 361 249
rect 395 215 429 249
rect 508 215 542 249
rect 630 215 664 249
rect 698 215 732 249
rect 806 215 840 249
rect 914 215 948 249
rect 1022 215 1056 249
rect 1090 215 1124 249
rect 1200 215 1234 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 96 485 162 527
rect 96 451 112 485
rect 146 451 162 485
rect 96 408 162 451
rect 96 374 112 408
rect 146 374 162 408
rect 196 477 232 493
rect 196 443 198 477
rect 196 386 232 443
rect 196 352 198 386
rect 268 485 334 527
rect 268 451 284 485
rect 318 451 334 485
rect 268 408 334 451
rect 268 374 284 408
rect 318 374 334 408
rect 368 477 406 493
rect 368 443 370 477
rect 404 443 406 477
rect 368 386 406 443
rect 440 481 506 527
rect 440 447 456 481
rect 490 447 506 481
rect 440 440 506 447
rect 540 477 612 493
rect 540 443 562 477
rect 596 443 612 477
rect 540 405 612 443
rect 657 489 723 527
rect 657 455 673 489
rect 707 455 723 489
rect 657 439 723 455
rect 757 477 824 493
rect 757 443 773 477
rect 807 443 824 477
rect 757 405 824 443
rect 858 489 911 527
rect 858 455 867 489
rect 901 455 911 489
rect 858 439 911 455
rect 1031 489 1097 493
rect 1031 455 1047 489
rect 1081 455 1097 489
rect 1031 421 1097 455
rect 1031 405 1047 421
rect 196 340 232 352
rect 368 352 370 386
rect 404 352 406 386
rect 368 340 406 352
rect 17 287 406 340
rect 440 387 1047 405
rect 1081 387 1097 421
rect 440 371 1097 387
rect 1203 485 1269 527
rect 1203 451 1219 485
rect 1253 451 1269 485
rect 1203 417 1269 451
rect 1203 383 1219 417
rect 1253 383 1269 417
rect 17 161 73 287
rect 440 253 474 371
rect 107 249 474 253
rect 107 215 123 249
rect 157 215 191 249
rect 225 215 259 249
rect 293 215 327 249
rect 361 215 395 249
rect 429 215 474 249
rect 107 213 474 215
rect 440 163 474 213
rect 508 289 856 337
rect 508 249 566 289
rect 542 215 566 249
rect 508 199 566 215
rect 611 249 748 255
rect 611 215 630 249
rect 664 215 698 249
rect 732 215 748 249
rect 611 207 748 215
rect 790 249 856 289
rect 790 215 806 249
rect 840 215 856 249
rect 790 207 856 215
rect 898 299 1258 337
rect 898 249 969 299
rect 898 215 914 249
rect 948 215 969 249
rect 898 207 969 215
rect 1006 249 1141 265
rect 1006 215 1022 249
rect 1056 215 1090 249
rect 1124 215 1141 249
rect 1006 207 1141 215
rect 1178 249 1258 299
rect 1178 215 1200 249
rect 1234 215 1258 249
rect 1178 207 1258 215
rect 834 169 1269 173
rect 17 127 321 161
rect 440 129 654 163
rect 688 129 704 163
rect 440 127 704 129
rect 834 135 850 169
rect 884 161 1269 169
rect 884 157 1219 161
rect 884 139 1047 157
rect 884 135 900 139
rect 119 123 321 127
rect 119 101 153 123
rect 19 59 35 93
rect 69 59 85 93
rect 19 17 85 59
rect 287 101 321 123
rect 119 51 153 67
rect 187 55 203 89
rect 237 55 253 89
rect 187 17 253 55
rect 834 101 900 135
rect 1031 123 1047 139
rect 1081 139 1219 157
rect 1081 123 1097 139
rect 834 93 850 101
rect 287 51 321 67
rect 355 59 371 93
rect 405 59 428 93
rect 355 17 428 59
rect 466 59 482 93
rect 516 67 850 93
rect 884 67 900 101
rect 516 59 900 67
rect 466 51 900 59
rect 934 89 997 105
rect 934 55 947 89
rect 981 55 997 89
rect 934 17 997 55
rect 1031 89 1097 123
rect 1203 127 1219 139
rect 1253 127 1269 161
rect 1031 55 1047 89
rect 1081 55 1097 89
rect 1031 51 1097 55
rect 1131 89 1169 105
rect 1131 55 1133 89
rect 1167 55 1169 89
rect 1131 17 1169 55
rect 1203 93 1269 127
rect 1203 59 1219 93
rect 1253 59 1269 93
rect 1203 51 1269 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel locali s 1224 289 1258 323 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 29 153 63 187 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 672 221 706 255 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 1040 221 1074 255 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 764 289 798 323 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o211a_4
rlabel metal1 s 0 -48 1288 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1288 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_END 770896
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 761900
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 6.440 0.000 
<< end >>
