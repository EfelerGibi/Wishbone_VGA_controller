magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 12 21 2016 203
rect 29 -17 63 21
<< locali >>
rect 1592 409 1650 493
rect 1232 357 1650 409
rect 1592 333 1650 357
rect 1768 333 1818 493
rect 1936 333 2007 493
rect 337 289 1146 323
rect 1592 289 2007 333
rect 337 255 371 289
rect 1112 255 1146 289
rect 98 215 371 255
rect 435 215 1078 255
rect 1112 215 1486 255
rect 1963 181 2007 289
rect 1676 129 2007 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 17 323 92 493
rect 126 367 176 527
rect 210 401 260 493
rect 294 435 344 527
rect 378 401 428 493
rect 462 435 512 527
rect 546 401 596 493
rect 630 435 680 527
rect 714 401 764 493
rect 210 357 764 401
rect 807 401 870 493
rect 904 435 954 527
rect 988 401 1038 493
rect 1072 435 1122 527
rect 1156 443 1550 493
rect 1156 401 1198 443
rect 807 357 1198 401
rect 1684 367 1734 527
rect 210 323 260 357
rect 1852 367 1902 527
rect 17 289 260 323
rect 1180 289 1554 323
rect 17 181 64 289
rect 1520 255 1554 289
rect 1520 215 1929 255
rect 17 129 352 181
rect 386 145 772 181
rect 386 95 436 145
rect 34 51 436 95
rect 470 17 504 111
rect 538 51 604 145
rect 638 17 672 111
rect 706 51 772 145
rect 807 17 862 181
rect 896 147 1642 181
rect 896 145 1486 147
rect 896 51 962 145
rect 996 17 1030 111
rect 1064 51 1130 145
rect 1164 17 1198 111
rect 1232 51 1298 145
rect 1332 17 1366 111
rect 1400 51 1466 145
rect 1500 17 1554 111
rect 1592 95 1642 147
rect 1592 61 1994 95
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< obsm1 >>
rect 201 320 259 329
rect 1213 320 1271 329
rect 201 292 1271 320
rect 201 283 259 292
rect 1213 283 1271 292
<< labels >>
rlabel locali s 435 215 1078 255 6 A
port 1 nsew signal input
rlabel locali s 1112 215 1486 255 6 B
port 2 nsew signal input
rlabel locali s 1112 255 1146 289 6 B
port 2 nsew signal input
rlabel locali s 98 215 371 255 6 B
port 2 nsew signal input
rlabel locali s 337 255 371 289 6 B
port 2 nsew signal input
rlabel locali s 337 289 1146 323 6 B
port 2 nsew signal input
rlabel metal1 s 0 -48 2024 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 12 21 2016 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 2062 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 2024 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 1676 129 2007 181 6 Y
port 7 nsew signal output
rlabel locali s 1963 181 2007 289 6 Y
port 7 nsew signal output
rlabel locali s 1592 289 2007 333 6 Y
port 7 nsew signal output
rlabel locali s 1936 333 2007 493 6 Y
port 7 nsew signal output
rlabel locali s 1768 333 1818 493 6 Y
port 7 nsew signal output
rlabel locali s 1592 333 1650 357 6 Y
port 7 nsew signal output
rlabel locali s 1232 357 1650 409 6 Y
port 7 nsew signal output
rlabel locali s 1592 409 1650 493 6 Y
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2024 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 610512
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 596472
<< end >>
