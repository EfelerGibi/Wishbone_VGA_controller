magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 404 157 588 203
rect 23 21 588 157
rect 29 -17 63 21
<< locali >>
rect 17 211 125 323
rect 514 299 627 493
rect 535 165 627 299
rect 514 51 627 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 401 97 493
rect 131 435 185 527
rect 231 427 285 493
rect 17 357 206 401
rect 159 265 206 357
rect 251 323 285 427
rect 323 401 375 493
rect 415 435 480 527
rect 323 357 480 401
rect 159 199 217 265
rect 251 211 406 323
rect 440 265 480 357
rect 159 177 206 199
rect 17 143 206 177
rect 17 51 97 143
rect 251 117 285 211
rect 440 199 501 265
rect 440 177 480 199
rect 131 17 185 109
rect 231 51 285 117
rect 323 143 480 177
rect 323 51 375 143
rect 415 17 480 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 17 211 125 323 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 23 21 588 157 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 404 157 588 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 514 51 627 165 6 X
port 6 nsew signal output
rlabel locali s 535 165 627 299 6 X
port 6 nsew signal output
rlabel locali s 514 299 627 493 6 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2903432
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2897572
<< end >>
