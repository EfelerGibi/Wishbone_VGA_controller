magic
tech sky130A
magscale 1 2
timestamp 1683767628
use sky130_fd_pr__hvdfl1sd__example_5595914180851  sky130_fd_pr__hvdfl1sd__example_5595914180851_0
timestamp 1683767628
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_5595914180851  sky130_fd_pr__hvdfl1sd__example_5595914180851_1
timestamp 1683767628
transform 1 0 800 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 15442750
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 15441888
<< end >>
