magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 505 157 712 203
rect 1195 157 1379 203
rect 1 21 1379 157
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 259 47 289 119
rect 364 47 394 119
rect 486 47 516 131
rect 604 47 634 177
rect 792 47 822 131
rect 876 47 906 131
rect 1064 47 1094 131
rect 1176 47 1206 131
rect 1271 47 1301 177
<< scpmoshvt >>
rect 79 369 109 497
rect 151 369 181 497
rect 256 413 286 497
rect 352 413 382 497
rect 470 413 500 497
rect 606 297 636 497
rect 792 303 822 431
rect 902 303 932 431
rect 1092 369 1122 497
rect 1176 369 1206 497
rect 1271 297 1301 497
<< ndiff >>
rect 27 103 79 131
rect 27 69 35 103
rect 69 69 79 103
rect 27 47 79 69
rect 109 89 163 131
rect 109 55 119 89
rect 153 55 163 89
rect 109 47 163 55
rect 193 119 244 131
rect 531 131 604 177
rect 436 119 486 131
rect 193 101 259 119
rect 193 67 203 101
rect 237 67 259 101
rect 193 47 259 67
rect 289 89 364 119
rect 289 55 309 89
rect 343 55 364 89
rect 289 47 364 55
rect 394 47 486 119
rect 516 119 604 131
rect 516 85 545 119
rect 579 85 604 119
rect 516 47 604 85
rect 634 101 686 177
rect 1221 131 1271 177
rect 634 67 644 101
rect 678 67 686 101
rect 634 47 686 67
rect 740 110 792 131
rect 740 76 748 110
rect 782 76 792 110
rect 740 47 792 76
rect 822 89 876 131
rect 822 55 832 89
rect 866 55 876 89
rect 822 47 876 55
rect 906 110 958 131
rect 906 76 916 110
rect 950 76 958 110
rect 906 47 958 76
rect 1012 109 1064 131
rect 1012 75 1020 109
rect 1054 75 1064 109
rect 1012 47 1064 75
rect 1094 47 1176 131
rect 1206 89 1271 131
rect 1206 55 1216 89
rect 1250 55 1271 89
rect 1206 47 1271 55
rect 1301 101 1353 177
rect 1301 67 1311 101
rect 1345 67 1353 101
rect 1301 47 1353 67
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 369 79 383
rect 109 369 151 497
rect 181 475 256 497
rect 181 441 201 475
rect 235 441 256 475
rect 181 413 256 441
rect 286 480 352 497
rect 286 446 302 480
rect 336 446 352 480
rect 286 413 352 446
rect 382 413 470 497
rect 500 489 606 497
rect 500 455 541 489
rect 575 455 606 489
rect 500 413 606 455
rect 181 369 241 413
rect 556 297 606 413
rect 636 477 688 497
rect 636 443 646 477
rect 680 443 688 477
rect 636 431 688 443
rect 837 485 887 497
rect 837 451 845 485
rect 879 451 887 485
rect 837 431 887 451
rect 1040 485 1092 497
rect 1040 451 1048 485
rect 1082 451 1092 485
rect 636 297 686 431
rect 742 361 792 431
rect 740 349 792 361
rect 740 315 748 349
rect 782 315 792 349
rect 740 303 792 315
rect 822 303 902 431
rect 932 349 984 431
rect 1040 369 1092 451
rect 1122 442 1176 497
rect 1122 408 1132 442
rect 1166 408 1176 442
rect 1122 369 1176 408
rect 1206 489 1271 497
rect 1206 455 1222 489
rect 1256 455 1271 489
rect 1206 369 1271 455
rect 932 315 942 349
rect 976 315 984 349
rect 932 303 984 315
rect 1221 297 1271 369
rect 1301 448 1353 497
rect 1301 414 1311 448
rect 1345 414 1353 448
rect 1301 380 1353 414
rect 1301 346 1311 380
rect 1345 346 1353 380
rect 1301 297 1353 346
<< ndiffc >>
rect 35 69 69 103
rect 119 55 153 89
rect 203 67 237 101
rect 309 55 343 89
rect 545 85 579 119
rect 644 67 678 101
rect 748 76 782 110
rect 832 55 866 89
rect 916 76 950 110
rect 1020 75 1054 109
rect 1216 55 1250 89
rect 1311 67 1345 101
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 201 441 235 475
rect 302 446 336 480
rect 541 455 575 489
rect 646 443 680 477
rect 845 451 879 485
rect 1048 451 1082 485
rect 748 315 782 349
rect 1132 408 1166 442
rect 1222 455 1256 489
rect 942 315 976 349
rect 1311 414 1345 448
rect 1311 346 1345 380
<< poly >>
rect 79 497 109 523
rect 151 497 181 523
rect 256 497 286 523
rect 352 497 382 523
rect 470 497 500 523
rect 606 497 636 523
rect 79 265 109 369
rect 21 249 109 265
rect 21 215 31 249
rect 65 215 109 249
rect 21 199 109 215
rect 151 265 181 369
rect 256 273 286 413
rect 352 381 382 413
rect 470 381 500 413
rect 328 365 382 381
rect 328 331 338 365
rect 372 331 382 365
rect 328 315 382 331
rect 464 365 518 381
rect 464 331 474 365
rect 508 331 518 365
rect 464 315 518 331
rect 151 249 214 265
rect 151 215 170 249
rect 204 215 214 249
rect 256 243 394 273
rect 151 199 214 215
rect 364 207 394 243
rect 79 131 109 199
rect 163 131 193 199
rect 256 191 322 201
rect 256 157 272 191
rect 306 157 322 191
rect 256 147 322 157
rect 364 191 418 207
rect 364 157 374 191
rect 408 157 418 191
rect 259 119 289 147
rect 364 141 418 157
rect 364 119 394 141
rect 486 131 516 315
rect 792 431 822 523
rect 902 431 932 523
rect 1092 497 1122 523
rect 1176 497 1206 523
rect 1271 497 1301 523
rect 1092 331 1122 369
rect 1056 321 1122 331
rect 606 265 636 297
rect 792 265 822 303
rect 902 265 932 303
rect 1056 287 1072 321
rect 1106 287 1122 321
rect 1056 277 1122 287
rect 558 249 636 265
rect 558 215 568 249
rect 602 215 636 249
rect 558 199 636 215
rect 784 255 850 265
rect 784 221 800 255
rect 834 221 850 255
rect 784 211 850 221
rect 902 249 986 265
rect 902 215 942 249
rect 976 215 986 249
rect 604 177 634 199
rect 792 131 822 211
rect 902 176 986 215
rect 876 146 986 176
rect 876 131 906 146
rect 1064 131 1094 277
rect 1176 237 1206 369
rect 1271 265 1301 297
rect 1136 227 1206 237
rect 1136 193 1152 227
rect 1186 193 1206 227
rect 1248 249 1302 265
rect 1248 215 1258 249
rect 1292 215 1302 249
rect 1248 199 1302 215
rect 1136 183 1206 193
rect 1176 131 1206 183
rect 1271 177 1301 199
rect 79 21 109 47
rect 163 21 193 47
rect 259 21 289 47
rect 364 21 394 47
rect 486 21 516 47
rect 604 21 634 47
rect 792 21 822 47
rect 876 21 906 47
rect 1064 21 1094 47
rect 1176 21 1206 47
rect 1271 21 1301 47
<< polycont >>
rect 31 215 65 249
rect 338 331 372 365
rect 474 331 508 365
rect 170 215 204 249
rect 272 157 306 191
rect 374 157 408 191
rect 1072 287 1106 321
rect 568 215 602 249
rect 800 221 834 255
rect 942 215 976 249
rect 1152 193 1186 227
rect 1258 215 1292 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 17 485 69 527
rect 17 451 35 485
rect 17 417 69 451
rect 17 383 35 417
rect 17 367 69 383
rect 108 475 251 493
rect 108 441 201 475
rect 235 441 251 475
rect 108 425 251 441
rect 285 480 440 493
rect 285 446 302 480
rect 336 446 440 480
rect 285 425 440 446
rect 108 351 142 425
rect 17 249 68 333
rect 17 215 31 249
rect 65 215 68 249
rect 17 191 68 215
rect 102 292 142 351
rect 102 157 136 292
rect 176 289 247 391
rect 281 365 372 391
rect 281 331 338 365
rect 281 323 372 331
rect 281 289 305 323
rect 339 289 372 323
rect 176 265 238 289
rect 281 265 372 289
rect 170 249 238 265
rect 204 215 238 249
rect 170 191 238 215
rect 272 241 372 265
rect 406 275 440 425
rect 474 489 602 527
rect 474 455 541 489
rect 575 455 602 489
rect 474 415 602 455
rect 636 477 680 493
rect 636 443 646 477
rect 716 485 1098 527
rect 716 451 845 485
rect 879 451 1048 485
rect 1082 451 1098 485
rect 636 417 680 443
rect 1132 442 1166 493
rect 1206 489 1272 527
rect 1206 455 1222 489
rect 1256 455 1272 489
rect 1206 451 1272 455
rect 636 383 1090 417
rect 636 381 680 383
rect 474 365 680 381
rect 508 331 680 365
rect 474 327 680 331
rect 474 315 508 327
rect 406 249 602 275
rect 406 241 568 249
rect 272 191 340 241
rect 465 215 568 241
rect 306 157 340 191
rect 17 123 238 157
rect 272 141 340 157
rect 374 191 431 207
rect 408 187 431 191
rect 374 153 397 157
rect 374 141 431 153
rect 465 199 602 215
rect 17 103 69 123
rect 17 69 35 103
rect 203 101 238 123
rect 465 107 499 199
rect 17 51 69 69
rect 103 55 119 89
rect 153 55 169 89
rect 103 17 169 55
rect 237 67 238 101
rect 203 51 238 67
rect 272 89 499 107
rect 272 55 309 89
rect 343 55 499 89
rect 272 51 499 55
rect 533 119 602 165
rect 533 85 545 119
rect 579 85 602 119
rect 533 17 602 85
rect 636 101 680 327
rect 636 67 644 101
rect 678 67 680 101
rect 636 51 680 67
rect 716 315 748 349
rect 782 315 798 349
rect 832 323 942 349
rect 716 187 750 315
rect 832 289 859 323
rect 893 315 942 323
rect 976 315 992 349
rect 893 299 992 315
rect 1028 321 1090 383
rect 1306 448 1363 493
rect 1166 408 1272 417
rect 1132 355 1272 408
rect 832 255 893 289
rect 1028 287 1072 321
rect 1106 287 1122 321
rect 1156 287 1272 355
rect 1306 414 1311 448
rect 1345 414 1363 448
rect 1306 380 1363 414
rect 1306 346 1311 380
rect 1345 346 1363 380
rect 1306 299 1363 346
rect 1238 265 1272 287
rect 784 221 800 255
rect 834 221 893 255
rect 716 153 767 187
rect 835 157 893 221
rect 942 253 986 265
rect 942 249 1202 253
rect 976 227 1202 249
rect 976 215 1152 227
rect 942 193 1152 215
rect 1186 193 1202 227
rect 942 191 1202 193
rect 1238 249 1292 265
rect 1238 215 1258 249
rect 1238 199 1292 215
rect 1238 157 1272 199
rect 1329 165 1363 299
rect 716 110 782 153
rect 835 123 966 157
rect 716 76 748 110
rect 916 110 966 123
rect 716 51 782 76
rect 816 55 832 89
rect 866 55 882 89
rect 816 17 882 55
rect 950 76 966 110
rect 916 51 966 76
rect 1002 123 1272 157
rect 1002 109 1054 123
rect 1002 75 1020 109
rect 1306 101 1363 165
rect 1002 51 1054 75
rect 1101 55 1216 89
rect 1250 55 1272 89
rect 1101 17 1272 55
rect 1306 67 1311 101
rect 1345 67 1363 101
rect 1306 51 1363 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 305 289 339 323
rect 397 157 408 187
rect 408 157 431 187
rect 397 153 431 157
rect 859 289 893 323
rect 767 153 801 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 293 323 351 329
rect 293 289 305 323
rect 339 320 351 323
rect 847 323 905 329
rect 847 320 859 323
rect 339 292 859 320
rect 339 289 351 292
rect 293 283 351 289
rect 847 289 859 292
rect 893 289 905 323
rect 847 283 905 289
rect 385 187 443 193
rect 385 153 397 187
rect 431 184 443 187
rect 755 187 813 193
rect 755 184 767 187
rect 431 156 767 184
rect 431 153 443 156
rect 385 147 443 153
rect 755 153 767 156
rect 801 153 813 187
rect 755 147 813 153
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 SCE
port 3 nsew signal input
flabel locali s 951 221 985 255 0 FreeSans 200 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1321 425 1355 459 0 FreeSans 200 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1321 357 1355 391 0 FreeSans 200 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 213 357 247 391 0 FreeSans 200 0 0 0 GATE
port 2 nsew signal input
flabel locali s 1321 85 1355 119 0 FreeSans 200 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 213 289 247 323 0 FreeSans 200 0 0 0 GATE
port 2 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 SCE
port 3 nsew signal input
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 sdlclkp_1
rlabel metal1 s 0 -48 1380 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1380 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1380 544
string GDS_END 419710
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 408734
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 6.900 0.000 
<< end >>
