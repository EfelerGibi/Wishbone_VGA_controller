magic
tech sky130A
magscale 1 2
timestamp 1683767628
use sky130_fd_pr__nfet_01v8__example_55959141808496  sky130_fd_pr__nfet_01v8__example_55959141808496_0
timestamp 1683767628
transform -1 0 1744 0 -1 358
box -1 0 417 1
use sky130_fd_pr__nfet_01v8__example_55959141808497  sky130_fd_pr__nfet_01v8__example_55959141808497_0
timestamp 1683767628
transform -1 0 1154 0 1 158
box -1 0 417 1
use sky130_fd_pr__nfet_01v8__example_55959141808498  sky130_fd_pr__nfet_01v8__example_55959141808498_0
timestamp 1683767628
transform -1 0 484 0 1 158
box -1 0 117 1
use sky130_fd_pr__nfet_01v8__example_55959141808498  sky130_fd_pr__nfet_01v8__example_55959141808498_1
timestamp 1683767628
transform -1 0 312 0 1 158
box -1 0 117 1
use sky130_fd_pr__nfet_01v8__example_55959141808582  sky130_fd_pr__nfet_01v8__example_55959141808582_0
timestamp 1683767628
transform -1 0 1186 0 -1 884
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808583  sky130_fd_pr__nfet_01v8__example_55959141808583_0
timestamp 1683767628
transform -1 0 438 0 -1 884
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808583  sky130_fd_pr__nfet_01v8__example_55959141808583_1
timestamp 1683767628
transform -1 0 750 0 -1 884
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808580  sky130_fd_pr__pfet_01v8__example_55959141808580_0
timestamp 1683767628
transform -1 0 1565 0 -1 964
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808580  sky130_fd_pr__pfet_01v8__example_55959141808580_1
timestamp 1683767628
transform 1 0 1621 0 -1 964
box -1 0 121 1
<< properties >>
string GDS_END 8119246
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8100062
<< end >>
