magic
tech sky130A
timestamp 1683767628
<< properties >>
string GDS_END 36672440
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 36671540
<< end >>
