magic
tech sky130B
timestamp 1683767628
<< properties >>
string GDS_END 4474770
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 4473934
<< end >>
