magic
tech sky130B
timestamp 1683767628
<< properties >>
string GDS_END 57392
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 57068
<< end >>
