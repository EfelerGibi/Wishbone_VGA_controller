magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 1 21 523 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 399 47 429 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 434 297 464 497
<< ndiff >>
rect 27 165 79 177
rect 27 131 35 165
rect 69 131 79 165
rect 27 97 79 131
rect 27 63 35 97
rect 69 63 79 97
rect 27 47 79 63
rect 109 165 163 177
rect 109 131 119 165
rect 153 131 163 165
rect 109 97 163 131
rect 109 63 119 97
rect 153 63 163 97
rect 109 47 163 63
rect 193 97 247 177
rect 193 63 203 97
rect 237 63 247 97
rect 193 47 247 63
rect 277 165 399 177
rect 277 131 290 165
rect 324 131 399 165
rect 277 97 399 131
rect 277 63 290 97
rect 324 63 399 97
rect 277 47 399 63
rect 429 165 497 177
rect 429 131 451 165
rect 485 131 497 165
rect 429 97 497 131
rect 429 63 451 97
rect 485 63 497 97
rect 429 47 497 63
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 297 163 497
rect 193 297 247 497
rect 277 477 434 497
rect 277 443 389 477
rect 423 443 434 477
rect 277 344 434 443
rect 277 310 389 344
rect 423 310 434 344
rect 277 297 434 310
rect 464 485 524 497
rect 464 451 482 485
rect 516 451 524 485
rect 464 417 524 451
rect 464 383 482 417
rect 516 383 524 417
rect 464 349 524 383
rect 464 315 482 349
rect 516 315 524 349
rect 464 297 524 315
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 119 131 153 165
rect 119 63 153 97
rect 203 63 237 97
rect 290 131 324 165
rect 290 63 324 97
rect 451 131 485 165
rect 451 63 485 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 389 443 423 477
rect 389 310 423 344
rect 482 451 516 485
rect 482 383 516 417
rect 482 315 516 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 434 497 464 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 434 265 464 297
rect 22 249 109 265
rect 22 215 34 249
rect 68 215 109 249
rect 22 199 109 215
rect 151 249 205 265
rect 151 215 161 249
rect 195 215 205 249
rect 151 199 205 215
rect 247 249 325 265
rect 247 215 275 249
rect 309 215 325 249
rect 247 199 325 215
rect 399 249 531 265
rect 399 215 485 249
rect 519 215 531 249
rect 399 199 531 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 399 177 429 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 399 21 429 47
<< polycont >>
rect 34 215 68 249
rect 161 215 195 249
rect 275 215 309 249
rect 485 215 519 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 18 485 88 527
rect 18 451 35 485
rect 69 451 88 485
rect 18 417 88 451
rect 18 383 35 417
rect 69 383 88 417
rect 18 349 88 383
rect 18 315 35 349
rect 69 315 88 349
rect 18 299 88 315
rect 18 249 88 265
rect 18 215 34 249
rect 68 215 88 249
rect 122 249 211 493
rect 292 265 340 481
rect 122 215 161 249
rect 195 215 211 249
rect 245 249 340 265
rect 245 215 275 249
rect 309 215 340 249
rect 389 477 432 493
rect 423 443 432 477
rect 389 344 432 443
rect 423 310 432 344
rect 35 165 69 181
rect 35 97 69 131
rect 35 17 69 63
rect 103 165 340 181
rect 103 131 119 165
rect 153 147 290 165
rect 153 131 169 147
rect 103 97 169 131
rect 274 131 290 147
rect 324 131 340 165
rect 103 63 119 97
rect 153 63 169 97
rect 103 51 169 63
rect 203 97 237 113
rect 203 17 237 63
rect 274 97 340 131
rect 274 63 290 97
rect 324 63 340 97
rect 274 51 340 63
rect 389 165 432 310
rect 466 485 535 527
rect 466 451 482 485
rect 516 451 535 485
rect 466 417 535 451
rect 466 383 482 417
rect 516 383 535 417
rect 466 349 535 383
rect 466 315 482 349
rect 516 315 535 349
rect 466 299 535 315
rect 466 249 535 265
rect 466 215 485 249
rect 519 215 535 249
rect 466 199 535 215
rect 389 131 451 165
rect 485 131 535 165
rect 389 97 535 131
rect 389 63 451 97
rect 485 63 535 97
rect 389 52 535 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
flabel locali s 398 85 432 119 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 122 289 156 323 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 398 153 432 187 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 487 221 521 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 490 85 524 119 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 122 425 156 459 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 122 357 156 391 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 398 221 432 255 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 398 289 432 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 398 357 432 391 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 398 425 432 459 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 o31ai_1
rlabel metal1 s 0 -48 552 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 552 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 552 544
string GDS_END 1430156
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1423882
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 2.760 0.000 
<< end >>
