magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 16 -26 72 30
<< locali >>
rect 0 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 17 440 1086 527
rect 334 126 402 292
rect 698 190 768 440
rect 17 17 1086 126
rect 0 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
rlabel metal1 s 0 -48 1104 48 8 VGND
port 1 nsew ground input
rlabel viali s 1041 -17 1075 17 8 VGND
port 1 nsew ground input
rlabel viali s 949 -17 983 17 8 VGND
port 1 nsew ground input
rlabel viali s 857 -17 891 17 8 VGND
port 1 nsew ground input
rlabel viali s 765 -17 799 17 8 VGND
port 1 nsew ground input
rlabel viali s 673 -17 707 17 8 VGND
port 1 nsew ground input
rlabel viali s 581 -17 615 17 8 VGND
port 1 nsew ground input
rlabel viali s 489 -17 523 17 8 VGND
port 1 nsew ground input
rlabel viali s 397 -17 431 17 8 VGND
port 1 nsew ground input
rlabel viali s 305 -17 339 17 8 VGND
port 1 nsew ground input
rlabel viali s 213 -17 247 17 8 VGND
port 1 nsew ground input
rlabel viali s 121 -17 155 17 8 VGND
port 1 nsew ground input
rlabel locali s 0 -17 1104 17 8 VGND
port 1 nsew ground input
rlabel locali s 17 17 1086 126 6 VGND
port 1 nsew ground input
rlabel locali s 334 126 402 292 6 VGND
port 1 nsew ground input
rlabel pwell s 16 -26 72 30 6 VNB
port 2 nsew ground input
rlabel nwell s -38 261 1142 582 6 VPB
port 3 nsew power input
rlabel metal1 s 0 496 1104 592 6 VPWR
port 4 nsew power input
rlabel viali s 1041 527 1075 561 6 VPWR
port 4 nsew power input
rlabel viali s 949 527 983 561 6 VPWR
port 4 nsew power input
rlabel viali s 857 527 891 561 6 VPWR
port 4 nsew power input
rlabel viali s 765 527 799 561 6 VPWR
port 4 nsew power input
rlabel viali s 673 527 707 561 6 VPWR
port 4 nsew power input
rlabel viali s 581 527 615 561 6 VPWR
port 4 nsew power input
rlabel viali s 489 527 523 561 6 VPWR
port 4 nsew power input
rlabel viali s 397 527 431 561 6 VPWR
port 4 nsew power input
rlabel viali s 305 527 339 561 6 VPWR
port 4 nsew power input
rlabel viali s 213 527 247 561 6 VPWR
port 4 nsew power input
rlabel viali s 121 527 155 561 6 VPWR
port 4 nsew power input
rlabel locali s 698 190 768 440 6 VPWR
port 4 nsew power input
rlabel locali s 17 440 1086 527 6 VPWR
port 4 nsew power input
rlabel locali s 0 527 1104 561 6 VPWR
port 4 nsew power input
<< properties >>
string FIXED_BBOX 0 0 1104 544
string LEFclass CORE SPACER
string LEFview TRUE
string GDS_END 3961718
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3957992
<< end >>
