magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< dnwell >>
tri -700 6714 -614 6800 se
rect -614 6714 764 6800
tri 764 6714 850 6800 sw
rect -700 -714 850 6714
tri -700 -800 -614 -714 ne
rect -614 -800 764 -714
tri 764 -800 850 -714 nw
<< nwell >>
rect -10 0 160 6000
<< pwell >>
rect -1166 7074 1316 7208
rect -1166 6026 -1032 7074
rect 1182 6026 1316 7074
rect -1166 -26 -574 6026
rect 724 -26 1316 6026
rect -1166 -1074 -1032 -26
rect 1182 -1074 1316 -26
rect -1166 -1208 1316 -1074
<< obsactive >>
rect -1240 -1282 1390 7282
<< locali >>
rect -1140 7158 1290 7182
rect -1140 7124 -988 7158
rect -954 7124 -916 7158
rect -882 7124 -844 7158
rect -810 7124 -772 7158
rect -738 7124 -700 7158
rect -666 7124 -628 7158
rect -594 7124 -556 7158
rect -522 7124 -484 7158
rect -450 7124 -412 7158
rect -378 7124 -340 7158
rect -306 7124 -268 7158
rect -234 7124 -196 7158
rect -162 7124 -124 7158
rect -90 7124 -52 7158
rect -18 7124 20 7158
rect 54 7124 92 7158
rect 126 7124 164 7158
rect 198 7124 236 7158
rect 270 7124 308 7158
rect 342 7124 380 7158
rect 414 7124 452 7158
rect 486 7124 524 7158
rect 558 7124 596 7158
rect 630 7124 668 7158
rect 702 7124 740 7158
rect 774 7124 812 7158
rect 846 7124 884 7158
rect 918 7124 956 7158
rect 990 7124 1028 7158
rect 1062 7124 1100 7158
rect 1134 7124 1290 7158
rect -1140 7100 1290 7124
rect -1140 7085 -1058 7100
rect -1140 7051 -1116 7085
rect -1082 7051 -1058 7085
rect -1140 7013 -1058 7051
rect -1140 6979 -1116 7013
rect -1082 6979 -1058 7013
rect -1140 6941 -1058 6979
rect -1140 6907 -1116 6941
rect -1082 6907 -1058 6941
rect -1140 6869 -1058 6907
rect -1140 6835 -1116 6869
rect -1082 6835 -1058 6869
rect -1140 6797 -1058 6835
rect -1140 6763 -1116 6797
rect -1082 6763 -1058 6797
rect -1140 6725 -1058 6763
rect -1140 6691 -1116 6725
rect -1082 6691 -1058 6725
rect -1140 6653 -1058 6691
rect -1140 6619 -1116 6653
rect -1082 6619 -1058 6653
rect -1140 6581 -1058 6619
rect -1140 6547 -1116 6581
rect -1082 6547 -1058 6581
rect -1140 6509 -1058 6547
rect -1140 6475 -1116 6509
rect -1082 6475 -1058 6509
rect -1140 6437 -1058 6475
rect -1140 6403 -1116 6437
rect -1082 6403 -1058 6437
rect -1140 6365 -1058 6403
rect -1140 6331 -1116 6365
rect -1082 6331 -1058 6365
rect -1140 6293 -1058 6331
rect -1140 6259 -1116 6293
rect -1082 6259 -1058 6293
rect -1140 6221 -1058 6259
rect -1140 6187 -1116 6221
rect -1082 6187 -1058 6221
rect -1140 6149 -1058 6187
rect -1140 6115 -1116 6149
rect -1082 6115 -1058 6149
rect -1140 6077 -1058 6115
rect -1140 6043 -1116 6077
rect -1082 6043 -1058 6077
rect -1140 6005 -1058 6043
rect -1140 5971 -1116 6005
rect -1082 5971 -1058 6005
rect 1208 7085 1290 7100
rect 1208 7051 1232 7085
rect 1266 7051 1290 7085
rect 1208 7013 1290 7051
rect 1208 6979 1232 7013
rect 1266 6979 1290 7013
rect 1208 6941 1290 6979
rect 1208 6907 1232 6941
rect 1266 6907 1290 6941
rect 1208 6869 1290 6907
rect 1208 6835 1232 6869
rect 1266 6835 1290 6869
rect 1208 6797 1290 6835
rect 1208 6763 1232 6797
rect 1266 6763 1290 6797
rect 1208 6725 1290 6763
rect 1208 6691 1232 6725
rect 1266 6691 1290 6725
rect 1208 6653 1290 6691
rect 1208 6619 1232 6653
rect 1266 6619 1290 6653
rect 1208 6581 1290 6619
rect 1208 6547 1232 6581
rect 1266 6547 1290 6581
rect 1208 6509 1290 6547
rect 1208 6475 1232 6509
rect 1266 6475 1290 6509
rect 1208 6437 1290 6475
rect 1208 6403 1232 6437
rect 1266 6403 1290 6437
rect 1208 6365 1290 6403
rect 1208 6331 1232 6365
rect 1266 6331 1290 6365
rect 1208 6293 1290 6331
rect 1208 6259 1232 6293
rect 1266 6259 1290 6293
rect 1208 6221 1290 6259
rect 1208 6187 1232 6221
rect 1266 6187 1290 6221
rect 1208 6149 1290 6187
rect 1208 6115 1232 6149
rect 1266 6115 1290 6149
rect 1208 6077 1290 6115
rect 1208 6043 1232 6077
rect 1266 6043 1290 6077
rect 1208 6005 1290 6043
rect -1140 5933 -1058 5971
rect -1140 5899 -1116 5933
rect -1082 5899 -1058 5933
rect -1140 5861 -1058 5899
rect -1140 5827 -1116 5861
rect -1082 5827 -1058 5861
rect -1140 5789 -1058 5827
rect -1140 5755 -1116 5789
rect -1082 5755 -1058 5789
rect -1140 5717 -1058 5755
rect -1140 5683 -1116 5717
rect -1082 5683 -1058 5717
rect -1140 5645 -1058 5683
rect -1140 5611 -1116 5645
rect -1082 5611 -1058 5645
rect -1140 5573 -1058 5611
rect -1140 5539 -1116 5573
rect -1082 5539 -1058 5573
rect -1140 5501 -1058 5539
rect -1140 5467 -1116 5501
rect -1082 5467 -1058 5501
rect -1140 5429 -1058 5467
rect -1140 5395 -1116 5429
rect -1082 5395 -1058 5429
rect -1140 5357 -1058 5395
rect -1140 5323 -1116 5357
rect -1082 5323 -1058 5357
rect -1140 5285 -1058 5323
rect -1140 5251 -1116 5285
rect -1082 5251 -1058 5285
rect -1140 5213 -1058 5251
rect -1140 5179 -1116 5213
rect -1082 5179 -1058 5213
rect -1140 5141 -1058 5179
rect -1140 5107 -1116 5141
rect -1082 5107 -1058 5141
rect -1140 5069 -1058 5107
rect -1140 5035 -1116 5069
rect -1082 5035 -1058 5069
rect -1140 4997 -1058 5035
rect -1140 4963 -1116 4997
rect -1082 4963 -1058 4997
rect -1140 4925 -1058 4963
rect -1140 4891 -1116 4925
rect -1082 4891 -1058 4925
rect -1140 4853 -1058 4891
rect -1140 4819 -1116 4853
rect -1082 4819 -1058 4853
rect -1140 4781 -1058 4819
rect -1140 4747 -1116 4781
rect -1082 4747 -1058 4781
rect -1140 4709 -1058 4747
rect -1140 4675 -1116 4709
rect -1082 4675 -1058 4709
rect -1140 4637 -1058 4675
rect -1140 4603 -1116 4637
rect -1082 4603 -1058 4637
rect -1140 4565 -1058 4603
rect -1140 4531 -1116 4565
rect -1082 4531 -1058 4565
rect -1140 4493 -1058 4531
rect -1140 4459 -1116 4493
rect -1082 4459 -1058 4493
rect -1140 4421 -1058 4459
rect -1140 4387 -1116 4421
rect -1082 4387 -1058 4421
rect -1140 4349 -1058 4387
rect -1140 4315 -1116 4349
rect -1082 4315 -1058 4349
rect -1140 4277 -1058 4315
rect -1140 4243 -1116 4277
rect -1082 4243 -1058 4277
rect -1140 4205 -1058 4243
rect -1140 4171 -1116 4205
rect -1082 4171 -1058 4205
rect -1140 4133 -1058 4171
rect -1140 4099 -1116 4133
rect -1082 4099 -1058 4133
rect -1140 4061 -1058 4099
rect -1140 4027 -1116 4061
rect -1082 4027 -1058 4061
rect -1140 3989 -1058 4027
rect -1140 3955 -1116 3989
rect -1082 3955 -1058 3989
rect -1140 3917 -1058 3955
rect -1140 3883 -1116 3917
rect -1082 3883 -1058 3917
rect -1140 3845 -1058 3883
rect -1140 3811 -1116 3845
rect -1082 3811 -1058 3845
rect -1140 3773 -1058 3811
rect -1140 3739 -1116 3773
rect -1082 3739 -1058 3773
rect -1140 3701 -1058 3739
rect -1140 3667 -1116 3701
rect -1082 3667 -1058 3701
rect -1140 3629 -1058 3667
rect -1140 3595 -1116 3629
rect -1082 3595 -1058 3629
rect -1140 3557 -1058 3595
rect -1140 3523 -1116 3557
rect -1082 3523 -1058 3557
rect -1140 3485 -1058 3523
rect -1140 3451 -1116 3485
rect -1082 3451 -1058 3485
rect -1140 3413 -1058 3451
rect -1140 3379 -1116 3413
rect -1082 3379 -1058 3413
rect -1140 3341 -1058 3379
rect -1140 3307 -1116 3341
rect -1082 3307 -1058 3341
rect -1140 3269 -1058 3307
rect -1140 3235 -1116 3269
rect -1082 3235 -1058 3269
rect -1140 3197 -1058 3235
rect -1140 3163 -1116 3197
rect -1082 3163 -1058 3197
rect -1140 3125 -1058 3163
rect -1140 3091 -1116 3125
rect -1082 3091 -1058 3125
rect -1140 3053 -1058 3091
rect -1140 3019 -1116 3053
rect -1082 3019 -1058 3053
rect -1140 2981 -1058 3019
rect -1140 2947 -1116 2981
rect -1082 2947 -1058 2981
rect -1140 2909 -1058 2947
rect -1140 2875 -1116 2909
rect -1082 2875 -1058 2909
rect -1140 2837 -1058 2875
rect -1140 2803 -1116 2837
rect -1082 2803 -1058 2837
rect -1140 2765 -1058 2803
rect -1140 2731 -1116 2765
rect -1082 2731 -1058 2765
rect -1140 2693 -1058 2731
rect -1140 2659 -1116 2693
rect -1082 2659 -1058 2693
rect -1140 2621 -1058 2659
rect -1140 2587 -1116 2621
rect -1082 2587 -1058 2621
rect -1140 2549 -1058 2587
rect -1140 2515 -1116 2549
rect -1082 2515 -1058 2549
rect -1140 2477 -1058 2515
rect -1140 2443 -1116 2477
rect -1082 2443 -1058 2477
rect -1140 2405 -1058 2443
rect -1140 2371 -1116 2405
rect -1082 2371 -1058 2405
rect -1140 2333 -1058 2371
rect -1140 2299 -1116 2333
rect -1082 2299 -1058 2333
rect -1140 2261 -1058 2299
rect -1140 2227 -1116 2261
rect -1082 2227 -1058 2261
rect -1140 2189 -1058 2227
rect -1140 2155 -1116 2189
rect -1082 2155 -1058 2189
rect -1140 2117 -1058 2155
rect -1140 2083 -1116 2117
rect -1082 2083 -1058 2117
rect -1140 2045 -1058 2083
rect -1140 2011 -1116 2045
rect -1082 2011 -1058 2045
rect -1140 1973 -1058 2011
rect -1140 1939 -1116 1973
rect -1082 1939 -1058 1973
rect -1140 1901 -1058 1939
rect -1140 1867 -1116 1901
rect -1082 1867 -1058 1901
rect -1140 1829 -1058 1867
rect -1140 1795 -1116 1829
rect -1082 1795 -1058 1829
rect -1140 1757 -1058 1795
rect -1140 1723 -1116 1757
rect -1082 1723 -1058 1757
rect -1140 1685 -1058 1723
rect -1140 1651 -1116 1685
rect -1082 1651 -1058 1685
rect -1140 1613 -1058 1651
rect -1140 1579 -1116 1613
rect -1082 1579 -1058 1613
rect -1140 1541 -1058 1579
rect -1140 1507 -1116 1541
rect -1082 1507 -1058 1541
rect -1140 1469 -1058 1507
rect -1140 1435 -1116 1469
rect -1082 1435 -1058 1469
rect -1140 1397 -1058 1435
rect -1140 1363 -1116 1397
rect -1082 1363 -1058 1397
rect -1140 1325 -1058 1363
rect -1140 1291 -1116 1325
rect -1082 1291 -1058 1325
rect -1140 1253 -1058 1291
rect -1140 1219 -1116 1253
rect -1082 1219 -1058 1253
rect -1140 1181 -1058 1219
rect -1140 1147 -1116 1181
rect -1082 1147 -1058 1181
rect -1140 1109 -1058 1147
rect -1140 1075 -1116 1109
rect -1082 1075 -1058 1109
rect -1140 1037 -1058 1075
rect -1140 1003 -1116 1037
rect -1082 1003 -1058 1037
rect -1140 965 -1058 1003
rect -1140 931 -1116 965
rect -1082 931 -1058 965
rect -1140 893 -1058 931
rect -1140 859 -1116 893
rect -1082 859 -1058 893
rect -1140 821 -1058 859
rect -1140 787 -1116 821
rect -1082 787 -1058 821
rect -1140 749 -1058 787
rect -1140 715 -1116 749
rect -1082 715 -1058 749
rect -1140 677 -1058 715
rect -1140 643 -1116 677
rect -1082 643 -1058 677
rect -1140 605 -1058 643
rect -1140 571 -1116 605
rect -1082 571 -1058 605
rect -1140 533 -1058 571
rect -1140 499 -1116 533
rect -1082 499 -1058 533
rect -1140 461 -1058 499
rect -1140 427 -1116 461
rect -1082 427 -1058 461
rect -1140 389 -1058 427
rect -1140 355 -1116 389
rect -1082 355 -1058 389
rect -1140 317 -1058 355
rect -1140 283 -1116 317
rect -1082 283 -1058 317
rect -1140 245 -1058 283
rect -1140 211 -1116 245
rect -1082 211 -1058 245
rect -1140 173 -1058 211
rect -1140 139 -1116 173
rect -1082 139 -1058 173
rect -1140 101 -1058 139
rect -1140 67 -1116 101
rect -1082 67 -1058 101
rect -1140 29 -1058 67
rect -1140 -5 -1116 29
rect -1082 -5 -1058 29
rect -962 5969 -896 5991
rect -962 5935 -946 5969
rect -912 5935 -896 5969
rect 1046 5969 1112 5991
rect -962 5897 -896 5935
rect -962 5863 -946 5897
rect -912 5863 -896 5897
rect -962 5825 -896 5863
rect -962 5791 -946 5825
rect -912 5791 -896 5825
rect -962 5753 -896 5791
rect -962 5719 -946 5753
rect -912 5719 -896 5753
rect -962 5681 -896 5719
rect -962 5647 -946 5681
rect -912 5647 -896 5681
rect -962 5609 -896 5647
rect -962 5575 -946 5609
rect -912 5575 -896 5609
rect -962 5537 -896 5575
rect -962 5503 -946 5537
rect -912 5503 -896 5537
rect -962 5465 -896 5503
rect -962 5431 -946 5465
rect -912 5431 -896 5465
rect -962 5393 -896 5431
rect -962 5359 -946 5393
rect -912 5359 -896 5393
rect -962 5321 -896 5359
rect -962 5287 -946 5321
rect -912 5287 -896 5321
rect -962 5249 -896 5287
rect -962 5215 -946 5249
rect -912 5215 -896 5249
rect -962 5177 -896 5215
rect -962 5143 -946 5177
rect -912 5143 -896 5177
rect -962 5105 -896 5143
rect -962 5071 -946 5105
rect -912 5071 -896 5105
rect -962 5033 -896 5071
rect -962 4999 -946 5033
rect -912 4999 -896 5033
rect -962 4961 -896 4999
rect -962 4927 -946 4961
rect -912 4927 -896 4961
rect -962 4889 -896 4927
rect -962 4855 -946 4889
rect -912 4855 -896 4889
rect -962 4817 -896 4855
rect -962 4783 -946 4817
rect -912 4783 -896 4817
rect -962 4745 -896 4783
rect -962 4711 -946 4745
rect -912 4711 -896 4745
rect -962 4673 -896 4711
rect -962 4639 -946 4673
rect -912 4639 -896 4673
rect -962 4601 -896 4639
rect -962 4567 -946 4601
rect -912 4567 -896 4601
rect -962 4529 -896 4567
rect -962 4495 -946 4529
rect -912 4495 -896 4529
rect -962 4457 -896 4495
rect -962 4423 -946 4457
rect -912 4423 -896 4457
rect -962 4385 -896 4423
rect -962 4351 -946 4385
rect -912 4351 -896 4385
rect -962 4313 -896 4351
rect -962 4279 -946 4313
rect -912 4279 -896 4313
rect -962 4241 -896 4279
rect -962 4207 -946 4241
rect -912 4207 -896 4241
rect -962 4169 -896 4207
rect -962 4135 -946 4169
rect -912 4135 -896 4169
rect -962 4097 -896 4135
rect -962 4063 -946 4097
rect -912 4063 -896 4097
rect -962 4025 -896 4063
rect -962 3991 -946 4025
rect -912 3991 -896 4025
rect -962 3953 -896 3991
rect -962 3919 -946 3953
rect -912 3919 -896 3953
rect -962 3881 -896 3919
rect -962 3847 -946 3881
rect -912 3847 -896 3881
rect -962 3809 -896 3847
rect -962 3775 -946 3809
rect -912 3775 -896 3809
rect -962 3737 -896 3775
rect -962 3703 -946 3737
rect -912 3703 -896 3737
rect -962 3665 -896 3703
rect -962 3631 -946 3665
rect -912 3631 -896 3665
rect -962 3593 -896 3631
rect -962 3559 -946 3593
rect -912 3559 -896 3593
rect -962 3521 -896 3559
rect -962 3487 -946 3521
rect -912 3487 -896 3521
rect -962 3449 -896 3487
rect -962 3415 -946 3449
rect -912 3415 -896 3449
rect -962 3377 -896 3415
rect -962 3343 -946 3377
rect -912 3343 -896 3377
rect -962 3305 -896 3343
rect -962 3271 -946 3305
rect -912 3271 -896 3305
rect -962 3233 -896 3271
rect -962 3199 -946 3233
rect -912 3199 -896 3233
rect -962 3161 -896 3199
rect -962 3127 -946 3161
rect -912 3127 -896 3161
rect -962 3089 -896 3127
rect -962 3055 -946 3089
rect -912 3055 -896 3089
rect -962 3017 -896 3055
rect -962 2983 -946 3017
rect -912 2983 -896 3017
rect -962 2945 -896 2983
rect -962 2911 -946 2945
rect -912 2911 -896 2945
rect -962 2873 -896 2911
rect -962 2839 -946 2873
rect -912 2839 -896 2873
rect -962 2801 -896 2839
rect -962 2767 -946 2801
rect -912 2767 -896 2801
rect -962 2729 -896 2767
rect -962 2695 -946 2729
rect -912 2695 -896 2729
rect -962 2657 -896 2695
rect -962 2623 -946 2657
rect -912 2623 -896 2657
rect -962 2585 -896 2623
rect -962 2551 -946 2585
rect -912 2551 -896 2585
rect -962 2513 -896 2551
rect -962 2479 -946 2513
rect -912 2479 -896 2513
rect -962 2441 -896 2479
rect -962 2407 -946 2441
rect -912 2407 -896 2441
rect -962 2369 -896 2407
rect -962 2335 -946 2369
rect -912 2335 -896 2369
rect -962 2297 -896 2335
rect -962 2263 -946 2297
rect -912 2263 -896 2297
rect -962 2225 -896 2263
rect -962 2191 -946 2225
rect -912 2191 -896 2225
rect -962 2153 -896 2191
rect -962 2119 -946 2153
rect -912 2119 -896 2153
rect -962 2081 -896 2119
rect -962 2047 -946 2081
rect -912 2047 -896 2081
rect -962 2009 -896 2047
rect -962 1975 -946 2009
rect -912 1975 -896 2009
rect -962 1937 -896 1975
rect -962 1903 -946 1937
rect -912 1903 -896 1937
rect -962 1865 -896 1903
rect -962 1831 -946 1865
rect -912 1831 -896 1865
rect -962 1793 -896 1831
rect -962 1759 -946 1793
rect -912 1759 -896 1793
rect -962 1721 -896 1759
rect -962 1687 -946 1721
rect -912 1687 -896 1721
rect -962 1649 -896 1687
rect -962 1615 -946 1649
rect -912 1615 -896 1649
rect -962 1577 -896 1615
rect -962 1543 -946 1577
rect -912 1543 -896 1577
rect -962 1505 -896 1543
rect -962 1471 -946 1505
rect -912 1471 -896 1505
rect -962 1433 -896 1471
rect -962 1399 -946 1433
rect -912 1399 -896 1433
rect -962 1361 -896 1399
rect -962 1327 -946 1361
rect -912 1327 -896 1361
rect -962 1289 -896 1327
rect -962 1255 -946 1289
rect -912 1255 -896 1289
rect -962 1217 -896 1255
rect -962 1183 -946 1217
rect -912 1183 -896 1217
rect -962 1145 -896 1183
rect -962 1111 -946 1145
rect -912 1111 -896 1145
rect -962 1073 -896 1111
rect -962 1039 -946 1073
rect -912 1039 -896 1073
rect -962 1001 -896 1039
rect -962 967 -946 1001
rect -912 967 -896 1001
rect -962 929 -896 967
rect -962 895 -946 929
rect -912 895 -896 929
rect -962 857 -896 895
rect -962 823 -946 857
rect -912 823 -896 857
rect -962 785 -896 823
rect -962 751 -946 785
rect -912 751 -896 785
rect -962 713 -896 751
rect -962 679 -946 713
rect -912 679 -896 713
rect -962 641 -896 679
rect -962 607 -946 641
rect -912 607 -896 641
rect -962 569 -896 607
rect -962 535 -946 569
rect -912 535 -896 569
rect -962 497 -896 535
rect -962 463 -946 497
rect -912 463 -896 497
rect -962 425 -896 463
rect -962 391 -946 425
rect -912 391 -896 425
rect -962 353 -896 391
rect -962 319 -946 353
rect -912 319 -896 353
rect -962 281 -896 319
rect -962 247 -946 281
rect -912 247 -896 281
rect -962 209 -896 247
rect -962 175 -946 209
rect -912 175 -896 209
rect -962 137 -896 175
rect -962 103 -946 137
rect -912 103 -896 137
rect -962 65 -896 103
rect -962 31 -946 65
rect -912 31 -896 65
rect 8 5933 142 5957
rect 8 67 22 5933
rect 128 67 142 5933
rect 8 43 142 67
rect 1046 5935 1062 5969
rect 1096 5935 1112 5969
rect 1046 5897 1112 5935
rect 1046 5863 1062 5897
rect 1096 5863 1112 5897
rect 1046 5825 1112 5863
rect 1046 5791 1062 5825
rect 1096 5791 1112 5825
rect 1046 5753 1112 5791
rect 1046 5719 1062 5753
rect 1096 5719 1112 5753
rect 1046 5681 1112 5719
rect 1046 5647 1062 5681
rect 1096 5647 1112 5681
rect 1046 5609 1112 5647
rect 1046 5575 1062 5609
rect 1096 5575 1112 5609
rect 1046 5537 1112 5575
rect 1046 5503 1062 5537
rect 1096 5503 1112 5537
rect 1046 5465 1112 5503
rect 1046 5431 1062 5465
rect 1096 5431 1112 5465
rect 1046 5393 1112 5431
rect 1046 5359 1062 5393
rect 1096 5359 1112 5393
rect 1046 5321 1112 5359
rect 1046 5287 1062 5321
rect 1096 5287 1112 5321
rect 1046 5249 1112 5287
rect 1046 5215 1062 5249
rect 1096 5215 1112 5249
rect 1046 5177 1112 5215
rect 1046 5143 1062 5177
rect 1096 5143 1112 5177
rect 1046 5105 1112 5143
rect 1046 5071 1062 5105
rect 1096 5071 1112 5105
rect 1046 5033 1112 5071
rect 1046 4999 1062 5033
rect 1096 4999 1112 5033
rect 1046 4961 1112 4999
rect 1046 4927 1062 4961
rect 1096 4927 1112 4961
rect 1046 4889 1112 4927
rect 1046 4855 1062 4889
rect 1096 4855 1112 4889
rect 1046 4817 1112 4855
rect 1046 4783 1062 4817
rect 1096 4783 1112 4817
rect 1046 4745 1112 4783
rect 1046 4711 1062 4745
rect 1096 4711 1112 4745
rect 1046 4673 1112 4711
rect 1046 4639 1062 4673
rect 1096 4639 1112 4673
rect 1046 4601 1112 4639
rect 1046 4567 1062 4601
rect 1096 4567 1112 4601
rect 1046 4529 1112 4567
rect 1046 4495 1062 4529
rect 1096 4495 1112 4529
rect 1046 4457 1112 4495
rect 1046 4423 1062 4457
rect 1096 4423 1112 4457
rect 1046 4385 1112 4423
rect 1046 4351 1062 4385
rect 1096 4351 1112 4385
rect 1046 4313 1112 4351
rect 1046 4279 1062 4313
rect 1096 4279 1112 4313
rect 1046 4241 1112 4279
rect 1046 4207 1062 4241
rect 1096 4207 1112 4241
rect 1046 4169 1112 4207
rect 1046 4135 1062 4169
rect 1096 4135 1112 4169
rect 1046 4097 1112 4135
rect 1046 4063 1062 4097
rect 1096 4063 1112 4097
rect 1046 4025 1112 4063
rect 1046 3991 1062 4025
rect 1096 3991 1112 4025
rect 1046 3953 1112 3991
rect 1046 3919 1062 3953
rect 1096 3919 1112 3953
rect 1046 3881 1112 3919
rect 1046 3847 1062 3881
rect 1096 3847 1112 3881
rect 1046 3809 1112 3847
rect 1046 3775 1062 3809
rect 1096 3775 1112 3809
rect 1046 3737 1112 3775
rect 1046 3703 1062 3737
rect 1096 3703 1112 3737
rect 1046 3665 1112 3703
rect 1046 3631 1062 3665
rect 1096 3631 1112 3665
rect 1046 3593 1112 3631
rect 1046 3559 1062 3593
rect 1096 3559 1112 3593
rect 1046 3521 1112 3559
rect 1046 3487 1062 3521
rect 1096 3487 1112 3521
rect 1046 3449 1112 3487
rect 1046 3415 1062 3449
rect 1096 3415 1112 3449
rect 1046 3377 1112 3415
rect 1046 3343 1062 3377
rect 1096 3343 1112 3377
rect 1046 3305 1112 3343
rect 1046 3271 1062 3305
rect 1096 3271 1112 3305
rect 1046 3233 1112 3271
rect 1046 3199 1062 3233
rect 1096 3199 1112 3233
rect 1046 3161 1112 3199
rect 1046 3127 1062 3161
rect 1096 3127 1112 3161
rect 1046 3089 1112 3127
rect 1046 3055 1062 3089
rect 1096 3055 1112 3089
rect 1046 3017 1112 3055
rect 1046 2983 1062 3017
rect 1096 2983 1112 3017
rect 1046 2945 1112 2983
rect 1046 2911 1062 2945
rect 1096 2911 1112 2945
rect 1046 2873 1112 2911
rect 1046 2839 1062 2873
rect 1096 2839 1112 2873
rect 1046 2801 1112 2839
rect 1046 2767 1062 2801
rect 1096 2767 1112 2801
rect 1046 2729 1112 2767
rect 1046 2695 1062 2729
rect 1096 2695 1112 2729
rect 1046 2657 1112 2695
rect 1046 2623 1062 2657
rect 1096 2623 1112 2657
rect 1046 2585 1112 2623
rect 1046 2551 1062 2585
rect 1096 2551 1112 2585
rect 1046 2513 1112 2551
rect 1046 2479 1062 2513
rect 1096 2479 1112 2513
rect 1046 2441 1112 2479
rect 1046 2407 1062 2441
rect 1096 2407 1112 2441
rect 1046 2369 1112 2407
rect 1046 2335 1062 2369
rect 1096 2335 1112 2369
rect 1046 2297 1112 2335
rect 1046 2263 1062 2297
rect 1096 2263 1112 2297
rect 1046 2225 1112 2263
rect 1046 2191 1062 2225
rect 1096 2191 1112 2225
rect 1046 2153 1112 2191
rect 1046 2119 1062 2153
rect 1096 2119 1112 2153
rect 1046 2081 1112 2119
rect 1046 2047 1062 2081
rect 1096 2047 1112 2081
rect 1046 2009 1112 2047
rect 1046 1975 1062 2009
rect 1096 1975 1112 2009
rect 1046 1937 1112 1975
rect 1046 1903 1062 1937
rect 1096 1903 1112 1937
rect 1046 1865 1112 1903
rect 1046 1831 1062 1865
rect 1096 1831 1112 1865
rect 1046 1793 1112 1831
rect 1046 1759 1062 1793
rect 1096 1759 1112 1793
rect 1046 1721 1112 1759
rect 1046 1687 1062 1721
rect 1096 1687 1112 1721
rect 1046 1649 1112 1687
rect 1046 1615 1062 1649
rect 1096 1615 1112 1649
rect 1046 1577 1112 1615
rect 1046 1543 1062 1577
rect 1096 1543 1112 1577
rect 1046 1505 1112 1543
rect 1046 1471 1062 1505
rect 1096 1471 1112 1505
rect 1046 1433 1112 1471
rect 1046 1399 1062 1433
rect 1096 1399 1112 1433
rect 1046 1361 1112 1399
rect 1046 1327 1062 1361
rect 1096 1327 1112 1361
rect 1046 1289 1112 1327
rect 1046 1255 1062 1289
rect 1096 1255 1112 1289
rect 1046 1217 1112 1255
rect 1046 1183 1062 1217
rect 1096 1183 1112 1217
rect 1046 1145 1112 1183
rect 1046 1111 1062 1145
rect 1096 1111 1112 1145
rect 1046 1073 1112 1111
rect 1046 1039 1062 1073
rect 1096 1039 1112 1073
rect 1046 1001 1112 1039
rect 1046 967 1062 1001
rect 1096 967 1112 1001
rect 1046 929 1112 967
rect 1046 895 1062 929
rect 1096 895 1112 929
rect 1046 857 1112 895
rect 1046 823 1062 857
rect 1096 823 1112 857
rect 1046 785 1112 823
rect 1046 751 1062 785
rect 1096 751 1112 785
rect 1046 713 1112 751
rect 1046 679 1062 713
rect 1096 679 1112 713
rect 1046 641 1112 679
rect 1046 607 1062 641
rect 1096 607 1112 641
rect 1046 569 1112 607
rect 1046 535 1062 569
rect 1096 535 1112 569
rect 1046 497 1112 535
rect 1046 463 1062 497
rect 1096 463 1112 497
rect 1046 425 1112 463
rect 1046 391 1062 425
rect 1096 391 1112 425
rect 1046 353 1112 391
rect 1046 319 1062 353
rect 1096 319 1112 353
rect 1046 281 1112 319
rect 1046 247 1062 281
rect 1096 247 1112 281
rect 1046 209 1112 247
rect 1046 175 1062 209
rect 1096 175 1112 209
rect 1046 137 1112 175
rect 1046 103 1062 137
rect 1096 103 1112 137
rect 1046 65 1112 103
rect -962 9 -896 31
rect 1046 31 1062 65
rect 1096 31 1112 65
rect 1046 9 1112 31
rect 1208 5971 1232 6005
rect 1266 5971 1290 6005
rect 1208 5933 1290 5971
rect 1208 5899 1232 5933
rect 1266 5899 1290 5933
rect 1208 5861 1290 5899
rect 1208 5827 1232 5861
rect 1266 5827 1290 5861
rect 1208 5789 1290 5827
rect 1208 5755 1232 5789
rect 1266 5755 1290 5789
rect 1208 5717 1290 5755
rect 1208 5683 1232 5717
rect 1266 5683 1290 5717
rect 1208 5645 1290 5683
rect 1208 5611 1232 5645
rect 1266 5611 1290 5645
rect 1208 5573 1290 5611
rect 1208 5539 1232 5573
rect 1266 5539 1290 5573
rect 1208 5501 1290 5539
rect 1208 5467 1232 5501
rect 1266 5467 1290 5501
rect 1208 5429 1290 5467
rect 1208 5395 1232 5429
rect 1266 5395 1290 5429
rect 1208 5357 1290 5395
rect 1208 5323 1232 5357
rect 1266 5323 1290 5357
rect 1208 5285 1290 5323
rect 1208 5251 1232 5285
rect 1266 5251 1290 5285
rect 1208 5213 1290 5251
rect 1208 5179 1232 5213
rect 1266 5179 1290 5213
rect 1208 5141 1290 5179
rect 1208 5107 1232 5141
rect 1266 5107 1290 5141
rect 1208 5069 1290 5107
rect 1208 5035 1232 5069
rect 1266 5035 1290 5069
rect 1208 4997 1290 5035
rect 1208 4963 1232 4997
rect 1266 4963 1290 4997
rect 1208 4925 1290 4963
rect 1208 4891 1232 4925
rect 1266 4891 1290 4925
rect 1208 4853 1290 4891
rect 1208 4819 1232 4853
rect 1266 4819 1290 4853
rect 1208 4781 1290 4819
rect 1208 4747 1232 4781
rect 1266 4747 1290 4781
rect 1208 4709 1290 4747
rect 1208 4675 1232 4709
rect 1266 4675 1290 4709
rect 1208 4637 1290 4675
rect 1208 4603 1232 4637
rect 1266 4603 1290 4637
rect 1208 4565 1290 4603
rect 1208 4531 1232 4565
rect 1266 4531 1290 4565
rect 1208 4493 1290 4531
rect 1208 4459 1232 4493
rect 1266 4459 1290 4493
rect 1208 4421 1290 4459
rect 1208 4387 1232 4421
rect 1266 4387 1290 4421
rect 1208 4349 1290 4387
rect 1208 4315 1232 4349
rect 1266 4315 1290 4349
rect 1208 4277 1290 4315
rect 1208 4243 1232 4277
rect 1266 4243 1290 4277
rect 1208 4205 1290 4243
rect 1208 4171 1232 4205
rect 1266 4171 1290 4205
rect 1208 4133 1290 4171
rect 1208 4099 1232 4133
rect 1266 4099 1290 4133
rect 1208 4061 1290 4099
rect 1208 4027 1232 4061
rect 1266 4027 1290 4061
rect 1208 3989 1290 4027
rect 1208 3955 1232 3989
rect 1266 3955 1290 3989
rect 1208 3917 1290 3955
rect 1208 3883 1232 3917
rect 1266 3883 1290 3917
rect 1208 3845 1290 3883
rect 1208 3811 1232 3845
rect 1266 3811 1290 3845
rect 1208 3773 1290 3811
rect 1208 3739 1232 3773
rect 1266 3739 1290 3773
rect 1208 3701 1290 3739
rect 1208 3667 1232 3701
rect 1266 3667 1290 3701
rect 1208 3629 1290 3667
rect 1208 3595 1232 3629
rect 1266 3595 1290 3629
rect 1208 3557 1290 3595
rect 1208 3523 1232 3557
rect 1266 3523 1290 3557
rect 1208 3485 1290 3523
rect 1208 3451 1232 3485
rect 1266 3451 1290 3485
rect 1208 3413 1290 3451
rect 1208 3379 1232 3413
rect 1266 3379 1290 3413
rect 1208 3341 1290 3379
rect 1208 3307 1232 3341
rect 1266 3307 1290 3341
rect 1208 3269 1290 3307
rect 1208 3235 1232 3269
rect 1266 3235 1290 3269
rect 1208 3197 1290 3235
rect 1208 3163 1232 3197
rect 1266 3163 1290 3197
rect 1208 3125 1290 3163
rect 1208 3091 1232 3125
rect 1266 3091 1290 3125
rect 1208 3053 1290 3091
rect 1208 3019 1232 3053
rect 1266 3019 1290 3053
rect 1208 2981 1290 3019
rect 1208 2947 1232 2981
rect 1266 2947 1290 2981
rect 1208 2909 1290 2947
rect 1208 2875 1232 2909
rect 1266 2875 1290 2909
rect 1208 2837 1290 2875
rect 1208 2803 1232 2837
rect 1266 2803 1290 2837
rect 1208 2765 1290 2803
rect 1208 2731 1232 2765
rect 1266 2731 1290 2765
rect 1208 2693 1290 2731
rect 1208 2659 1232 2693
rect 1266 2659 1290 2693
rect 1208 2621 1290 2659
rect 1208 2587 1232 2621
rect 1266 2587 1290 2621
rect 1208 2549 1290 2587
rect 1208 2515 1232 2549
rect 1266 2515 1290 2549
rect 1208 2477 1290 2515
rect 1208 2443 1232 2477
rect 1266 2443 1290 2477
rect 1208 2405 1290 2443
rect 1208 2371 1232 2405
rect 1266 2371 1290 2405
rect 1208 2333 1290 2371
rect 1208 2299 1232 2333
rect 1266 2299 1290 2333
rect 1208 2261 1290 2299
rect 1208 2227 1232 2261
rect 1266 2227 1290 2261
rect 1208 2189 1290 2227
rect 1208 2155 1232 2189
rect 1266 2155 1290 2189
rect 1208 2117 1290 2155
rect 1208 2083 1232 2117
rect 1266 2083 1290 2117
rect 1208 2045 1290 2083
rect 1208 2011 1232 2045
rect 1266 2011 1290 2045
rect 1208 1973 1290 2011
rect 1208 1939 1232 1973
rect 1266 1939 1290 1973
rect 1208 1901 1290 1939
rect 1208 1867 1232 1901
rect 1266 1867 1290 1901
rect 1208 1829 1290 1867
rect 1208 1795 1232 1829
rect 1266 1795 1290 1829
rect 1208 1757 1290 1795
rect 1208 1723 1232 1757
rect 1266 1723 1290 1757
rect 1208 1685 1290 1723
rect 1208 1651 1232 1685
rect 1266 1651 1290 1685
rect 1208 1613 1290 1651
rect 1208 1579 1232 1613
rect 1266 1579 1290 1613
rect 1208 1541 1290 1579
rect 1208 1507 1232 1541
rect 1266 1507 1290 1541
rect 1208 1469 1290 1507
rect 1208 1435 1232 1469
rect 1266 1435 1290 1469
rect 1208 1397 1290 1435
rect 1208 1363 1232 1397
rect 1266 1363 1290 1397
rect 1208 1325 1290 1363
rect 1208 1291 1232 1325
rect 1266 1291 1290 1325
rect 1208 1253 1290 1291
rect 1208 1219 1232 1253
rect 1266 1219 1290 1253
rect 1208 1181 1290 1219
rect 1208 1147 1232 1181
rect 1266 1147 1290 1181
rect 1208 1109 1290 1147
rect 1208 1075 1232 1109
rect 1266 1075 1290 1109
rect 1208 1037 1290 1075
rect 1208 1003 1232 1037
rect 1266 1003 1290 1037
rect 1208 965 1290 1003
rect 1208 931 1232 965
rect 1266 931 1290 965
rect 1208 893 1290 931
rect 1208 859 1232 893
rect 1266 859 1290 893
rect 1208 821 1290 859
rect 1208 787 1232 821
rect 1266 787 1290 821
rect 1208 749 1290 787
rect 1208 715 1232 749
rect 1266 715 1290 749
rect 1208 677 1290 715
rect 1208 643 1232 677
rect 1266 643 1290 677
rect 1208 605 1290 643
rect 1208 571 1232 605
rect 1266 571 1290 605
rect 1208 533 1290 571
rect 1208 499 1232 533
rect 1266 499 1290 533
rect 1208 461 1290 499
rect 1208 427 1232 461
rect 1266 427 1290 461
rect 1208 389 1290 427
rect 1208 355 1232 389
rect 1266 355 1290 389
rect 1208 317 1290 355
rect 1208 283 1232 317
rect 1266 283 1290 317
rect 1208 245 1290 283
rect 1208 211 1232 245
rect 1266 211 1290 245
rect 1208 173 1290 211
rect 1208 139 1232 173
rect 1266 139 1290 173
rect 1208 101 1290 139
rect 1208 67 1232 101
rect 1266 67 1290 101
rect 1208 29 1290 67
rect -1140 -43 -1058 -5
rect -1140 -77 -1116 -43
rect -1082 -77 -1058 -43
rect -1140 -115 -1058 -77
rect -1140 -149 -1116 -115
rect -1082 -149 -1058 -115
rect -1140 -187 -1058 -149
rect -1140 -221 -1116 -187
rect -1082 -221 -1058 -187
rect -1140 -259 -1058 -221
rect -1140 -293 -1116 -259
rect -1082 -293 -1058 -259
rect -1140 -331 -1058 -293
rect -1140 -365 -1116 -331
rect -1082 -365 -1058 -331
rect -1140 -403 -1058 -365
rect -1140 -437 -1116 -403
rect -1082 -437 -1058 -403
rect -1140 -475 -1058 -437
rect -1140 -509 -1116 -475
rect -1082 -509 -1058 -475
rect -1140 -547 -1058 -509
rect -1140 -581 -1116 -547
rect -1082 -581 -1058 -547
rect -1140 -619 -1058 -581
rect -1140 -653 -1116 -619
rect -1082 -653 -1058 -619
rect 1208 -5 1232 29
rect 1266 -5 1290 29
rect 1208 -43 1290 -5
rect 1208 -77 1232 -43
rect 1266 -77 1290 -43
rect 1208 -115 1290 -77
rect 1208 -149 1232 -115
rect 1266 -149 1290 -115
rect 1208 -187 1290 -149
rect 1208 -221 1232 -187
rect 1266 -221 1290 -187
rect 1208 -259 1290 -221
rect 1208 -293 1232 -259
rect 1266 -293 1290 -259
rect 1208 -331 1290 -293
rect 1208 -365 1232 -331
rect 1266 -365 1290 -331
rect 1208 -403 1290 -365
rect 1208 -437 1232 -403
rect 1266 -437 1290 -403
rect 1208 -475 1290 -437
rect 1208 -509 1232 -475
rect 1266 -509 1290 -475
rect 1208 -547 1290 -509
rect 1208 -581 1232 -547
rect 1266 -581 1290 -547
rect 1208 -619 1290 -581
rect -1140 -691 -1058 -653
rect -1140 -725 -1116 -691
rect -1082 -725 -1058 -691
rect -1140 -763 -1058 -725
rect -1140 -797 -1116 -763
rect -1082 -797 -1058 -763
rect -1140 -835 -1058 -797
rect -1140 -869 -1116 -835
rect -1082 -869 -1058 -835
rect -296 -659 460 -643
rect -296 -693 -280 -659
rect -246 -693 -206 -659
rect -172 -693 -132 -659
rect -98 -693 -58 -659
rect -24 -693 16 -659
rect 50 -693 90 -659
rect 124 -693 164 -659
rect 198 -693 238 -659
rect 272 -693 312 -659
rect 346 -693 386 -659
rect 420 -693 460 -659
rect -296 -733 460 -693
rect -296 -767 -280 -733
rect -246 -767 -206 -733
rect -172 -767 -132 -733
rect -98 -767 -58 -733
rect -24 -767 16 -733
rect 50 -767 90 -733
rect 124 -767 164 -733
rect 198 -767 238 -733
rect 272 -767 312 -733
rect 346 -767 386 -733
rect 420 -767 460 -733
rect -296 -807 460 -767
rect -296 -841 -280 -807
rect -246 -841 -206 -807
rect -172 -841 -132 -807
rect -98 -841 -58 -807
rect -24 -841 16 -807
rect 50 -841 90 -807
rect 124 -841 164 -807
rect 198 -841 238 -807
rect 272 -841 312 -807
rect 346 -841 386 -807
rect 420 -841 460 -807
rect -296 -857 460 -841
rect 1208 -653 1232 -619
rect 1266 -653 1290 -619
rect 1208 -691 1290 -653
rect 1208 -725 1232 -691
rect 1266 -725 1290 -691
rect 1208 -763 1290 -725
rect 1208 -797 1232 -763
rect 1266 -797 1290 -763
rect 1208 -835 1290 -797
rect -1140 -907 -1058 -869
rect -1140 -941 -1116 -907
rect -1082 -941 -1058 -907
rect -1140 -979 -1058 -941
rect -1140 -1013 -1116 -979
rect -1082 -1013 -1058 -979
rect -1140 -1051 -1058 -1013
rect -1140 -1085 -1116 -1051
rect -1082 -1085 -1058 -1051
rect -1140 -1100 -1058 -1085
rect 1208 -869 1232 -835
rect 1266 -869 1290 -835
rect 1208 -907 1290 -869
rect 1208 -941 1232 -907
rect 1266 -941 1290 -907
rect 1208 -979 1290 -941
rect 1208 -1013 1232 -979
rect 1266 -1013 1290 -979
rect 1208 -1051 1290 -1013
rect 1208 -1085 1232 -1051
rect 1266 -1085 1290 -1051
rect 1208 -1100 1290 -1085
rect -1140 -1124 1290 -1100
rect -1140 -1158 -988 -1124
rect -954 -1158 -916 -1124
rect -882 -1158 -844 -1124
rect -810 -1158 -772 -1124
rect -738 -1158 -700 -1124
rect -666 -1158 -628 -1124
rect -594 -1158 -556 -1124
rect -522 -1158 -484 -1124
rect -450 -1158 -412 -1124
rect -378 -1158 -340 -1124
rect -306 -1158 -268 -1124
rect -234 -1158 -196 -1124
rect -162 -1158 -124 -1124
rect -90 -1158 -52 -1124
rect -18 -1158 20 -1124
rect 54 -1158 92 -1124
rect 126 -1158 164 -1124
rect 198 -1158 236 -1124
rect 270 -1158 308 -1124
rect 342 -1158 380 -1124
rect 414 -1158 452 -1124
rect 486 -1158 524 -1124
rect 558 -1158 596 -1124
rect 630 -1158 668 -1124
rect 702 -1158 740 -1124
rect 774 -1158 812 -1124
rect 846 -1158 884 -1124
rect 918 -1158 956 -1124
rect 990 -1158 1028 -1124
rect 1062 -1158 1100 -1124
rect 1134 -1158 1290 -1124
rect -1140 -1182 1290 -1158
<< viali >>
rect -988 7124 -954 7158
rect -916 7124 -882 7158
rect -844 7124 -810 7158
rect -772 7124 -738 7158
rect -700 7124 -666 7158
rect -628 7124 -594 7158
rect -556 7124 -522 7158
rect -484 7124 -450 7158
rect -412 7124 -378 7158
rect -340 7124 -306 7158
rect -268 7124 -234 7158
rect -196 7124 -162 7158
rect -124 7124 -90 7158
rect -52 7124 -18 7158
rect 20 7124 54 7158
rect 92 7124 126 7158
rect 164 7124 198 7158
rect 236 7124 270 7158
rect 308 7124 342 7158
rect 380 7124 414 7158
rect 452 7124 486 7158
rect 524 7124 558 7158
rect 596 7124 630 7158
rect 668 7124 702 7158
rect 740 7124 774 7158
rect 812 7124 846 7158
rect 884 7124 918 7158
rect 956 7124 990 7158
rect 1028 7124 1062 7158
rect 1100 7124 1134 7158
rect -1116 7051 -1082 7085
rect -1116 6979 -1082 7013
rect -1116 6907 -1082 6941
rect -1116 6835 -1082 6869
rect -1116 6763 -1082 6797
rect -1116 6691 -1082 6725
rect -1116 6619 -1082 6653
rect -1116 6547 -1082 6581
rect -1116 6475 -1082 6509
rect -1116 6403 -1082 6437
rect -1116 6331 -1082 6365
rect -1116 6259 -1082 6293
rect -1116 6187 -1082 6221
rect -1116 6115 -1082 6149
rect -1116 6043 -1082 6077
rect -1116 5971 -1082 6005
rect 1232 7051 1266 7085
rect 1232 6979 1266 7013
rect 1232 6907 1266 6941
rect 1232 6835 1266 6869
rect 1232 6763 1266 6797
rect 1232 6691 1266 6725
rect 1232 6619 1266 6653
rect 1232 6547 1266 6581
rect 1232 6475 1266 6509
rect 1232 6403 1266 6437
rect 1232 6331 1266 6365
rect 1232 6259 1266 6293
rect 1232 6187 1266 6221
rect 1232 6115 1266 6149
rect 1232 6043 1266 6077
rect -1116 5899 -1082 5933
rect -1116 5827 -1082 5861
rect -1116 5755 -1082 5789
rect -1116 5683 -1082 5717
rect -1116 5611 -1082 5645
rect -1116 5539 -1082 5573
rect -1116 5467 -1082 5501
rect -1116 5395 -1082 5429
rect -1116 5323 -1082 5357
rect -1116 5251 -1082 5285
rect -1116 5179 -1082 5213
rect -1116 5107 -1082 5141
rect -1116 5035 -1082 5069
rect -1116 4963 -1082 4997
rect -1116 4891 -1082 4925
rect -1116 4819 -1082 4853
rect -1116 4747 -1082 4781
rect -1116 4675 -1082 4709
rect -1116 4603 -1082 4637
rect -1116 4531 -1082 4565
rect -1116 4459 -1082 4493
rect -1116 4387 -1082 4421
rect -1116 4315 -1082 4349
rect -1116 4243 -1082 4277
rect -1116 4171 -1082 4205
rect -1116 4099 -1082 4133
rect -1116 4027 -1082 4061
rect -1116 3955 -1082 3989
rect -1116 3883 -1082 3917
rect -1116 3811 -1082 3845
rect -1116 3739 -1082 3773
rect -1116 3667 -1082 3701
rect -1116 3595 -1082 3629
rect -1116 3523 -1082 3557
rect -1116 3451 -1082 3485
rect -1116 3379 -1082 3413
rect -1116 3307 -1082 3341
rect -1116 3235 -1082 3269
rect -1116 3163 -1082 3197
rect -1116 3091 -1082 3125
rect -1116 3019 -1082 3053
rect -1116 2947 -1082 2981
rect -1116 2875 -1082 2909
rect -1116 2803 -1082 2837
rect -1116 2731 -1082 2765
rect -1116 2659 -1082 2693
rect -1116 2587 -1082 2621
rect -1116 2515 -1082 2549
rect -1116 2443 -1082 2477
rect -1116 2371 -1082 2405
rect -1116 2299 -1082 2333
rect -1116 2227 -1082 2261
rect -1116 2155 -1082 2189
rect -1116 2083 -1082 2117
rect -1116 2011 -1082 2045
rect -1116 1939 -1082 1973
rect -1116 1867 -1082 1901
rect -1116 1795 -1082 1829
rect -1116 1723 -1082 1757
rect -1116 1651 -1082 1685
rect -1116 1579 -1082 1613
rect -1116 1507 -1082 1541
rect -1116 1435 -1082 1469
rect -1116 1363 -1082 1397
rect -1116 1291 -1082 1325
rect -1116 1219 -1082 1253
rect -1116 1147 -1082 1181
rect -1116 1075 -1082 1109
rect -1116 1003 -1082 1037
rect -1116 931 -1082 965
rect -1116 859 -1082 893
rect -1116 787 -1082 821
rect -1116 715 -1082 749
rect -1116 643 -1082 677
rect -1116 571 -1082 605
rect -1116 499 -1082 533
rect -1116 427 -1082 461
rect -1116 355 -1082 389
rect -1116 283 -1082 317
rect -1116 211 -1082 245
rect -1116 139 -1082 173
rect -1116 67 -1082 101
rect -1116 -5 -1082 29
rect -946 5935 -912 5969
rect -946 5863 -912 5897
rect -946 5791 -912 5825
rect -946 5719 -912 5753
rect -946 5647 -912 5681
rect -946 5575 -912 5609
rect -946 5503 -912 5537
rect -946 5431 -912 5465
rect -946 5359 -912 5393
rect -946 5287 -912 5321
rect -946 5215 -912 5249
rect -946 5143 -912 5177
rect -946 5071 -912 5105
rect -946 4999 -912 5033
rect -946 4927 -912 4961
rect -946 4855 -912 4889
rect -946 4783 -912 4817
rect -946 4711 -912 4745
rect -946 4639 -912 4673
rect -946 4567 -912 4601
rect -946 4495 -912 4529
rect -946 4423 -912 4457
rect -946 4351 -912 4385
rect -946 4279 -912 4313
rect -946 4207 -912 4241
rect -946 4135 -912 4169
rect -946 4063 -912 4097
rect -946 3991 -912 4025
rect -946 3919 -912 3953
rect -946 3847 -912 3881
rect -946 3775 -912 3809
rect -946 3703 -912 3737
rect -946 3631 -912 3665
rect -946 3559 -912 3593
rect -946 3487 -912 3521
rect -946 3415 -912 3449
rect -946 3343 -912 3377
rect -946 3271 -912 3305
rect -946 3199 -912 3233
rect -946 3127 -912 3161
rect -946 3055 -912 3089
rect -946 2983 -912 3017
rect -946 2911 -912 2945
rect -946 2839 -912 2873
rect -946 2767 -912 2801
rect -946 2695 -912 2729
rect -946 2623 -912 2657
rect -946 2551 -912 2585
rect -946 2479 -912 2513
rect -946 2407 -912 2441
rect -946 2335 -912 2369
rect -946 2263 -912 2297
rect -946 2191 -912 2225
rect -946 2119 -912 2153
rect -946 2047 -912 2081
rect -946 1975 -912 2009
rect -946 1903 -912 1937
rect -946 1831 -912 1865
rect -946 1759 -912 1793
rect -946 1687 -912 1721
rect -946 1615 -912 1649
rect -946 1543 -912 1577
rect -946 1471 -912 1505
rect -946 1399 -912 1433
rect -946 1327 -912 1361
rect -946 1255 -912 1289
rect -946 1183 -912 1217
rect -946 1111 -912 1145
rect -946 1039 -912 1073
rect -946 967 -912 1001
rect -946 895 -912 929
rect -946 823 -912 857
rect -946 751 -912 785
rect -946 679 -912 713
rect -946 607 -912 641
rect -946 535 -912 569
rect -946 463 -912 497
rect -946 391 -912 425
rect -946 319 -912 353
rect -946 247 -912 281
rect -946 175 -912 209
rect -946 103 -912 137
rect -946 31 -912 65
rect 22 67 128 5933
rect 1062 5935 1096 5969
rect 1062 5863 1096 5897
rect 1062 5791 1096 5825
rect 1062 5719 1096 5753
rect 1062 5647 1096 5681
rect 1062 5575 1096 5609
rect 1062 5503 1096 5537
rect 1062 5431 1096 5465
rect 1062 5359 1096 5393
rect 1062 5287 1096 5321
rect 1062 5215 1096 5249
rect 1062 5143 1096 5177
rect 1062 5071 1096 5105
rect 1062 4999 1096 5033
rect 1062 4927 1096 4961
rect 1062 4855 1096 4889
rect 1062 4783 1096 4817
rect 1062 4711 1096 4745
rect 1062 4639 1096 4673
rect 1062 4567 1096 4601
rect 1062 4495 1096 4529
rect 1062 4423 1096 4457
rect 1062 4351 1096 4385
rect 1062 4279 1096 4313
rect 1062 4207 1096 4241
rect 1062 4135 1096 4169
rect 1062 4063 1096 4097
rect 1062 3991 1096 4025
rect 1062 3919 1096 3953
rect 1062 3847 1096 3881
rect 1062 3775 1096 3809
rect 1062 3703 1096 3737
rect 1062 3631 1096 3665
rect 1062 3559 1096 3593
rect 1062 3487 1096 3521
rect 1062 3415 1096 3449
rect 1062 3343 1096 3377
rect 1062 3271 1096 3305
rect 1062 3199 1096 3233
rect 1062 3127 1096 3161
rect 1062 3055 1096 3089
rect 1062 2983 1096 3017
rect 1062 2911 1096 2945
rect 1062 2839 1096 2873
rect 1062 2767 1096 2801
rect 1062 2695 1096 2729
rect 1062 2623 1096 2657
rect 1062 2551 1096 2585
rect 1062 2479 1096 2513
rect 1062 2407 1096 2441
rect 1062 2335 1096 2369
rect 1062 2263 1096 2297
rect 1062 2191 1096 2225
rect 1062 2119 1096 2153
rect 1062 2047 1096 2081
rect 1062 1975 1096 2009
rect 1062 1903 1096 1937
rect 1062 1831 1096 1865
rect 1062 1759 1096 1793
rect 1062 1687 1096 1721
rect 1062 1615 1096 1649
rect 1062 1543 1096 1577
rect 1062 1471 1096 1505
rect 1062 1399 1096 1433
rect 1062 1327 1096 1361
rect 1062 1255 1096 1289
rect 1062 1183 1096 1217
rect 1062 1111 1096 1145
rect 1062 1039 1096 1073
rect 1062 967 1096 1001
rect 1062 895 1096 929
rect 1062 823 1096 857
rect 1062 751 1096 785
rect 1062 679 1096 713
rect 1062 607 1096 641
rect 1062 535 1096 569
rect 1062 463 1096 497
rect 1062 391 1096 425
rect 1062 319 1096 353
rect 1062 247 1096 281
rect 1062 175 1096 209
rect 1062 103 1096 137
rect 1062 31 1096 65
rect 1232 5971 1266 6005
rect 1232 5899 1266 5933
rect 1232 5827 1266 5861
rect 1232 5755 1266 5789
rect 1232 5683 1266 5717
rect 1232 5611 1266 5645
rect 1232 5539 1266 5573
rect 1232 5467 1266 5501
rect 1232 5395 1266 5429
rect 1232 5323 1266 5357
rect 1232 5251 1266 5285
rect 1232 5179 1266 5213
rect 1232 5107 1266 5141
rect 1232 5035 1266 5069
rect 1232 4963 1266 4997
rect 1232 4891 1266 4925
rect 1232 4819 1266 4853
rect 1232 4747 1266 4781
rect 1232 4675 1266 4709
rect 1232 4603 1266 4637
rect 1232 4531 1266 4565
rect 1232 4459 1266 4493
rect 1232 4387 1266 4421
rect 1232 4315 1266 4349
rect 1232 4243 1266 4277
rect 1232 4171 1266 4205
rect 1232 4099 1266 4133
rect 1232 4027 1266 4061
rect 1232 3955 1266 3989
rect 1232 3883 1266 3917
rect 1232 3811 1266 3845
rect 1232 3739 1266 3773
rect 1232 3667 1266 3701
rect 1232 3595 1266 3629
rect 1232 3523 1266 3557
rect 1232 3451 1266 3485
rect 1232 3379 1266 3413
rect 1232 3307 1266 3341
rect 1232 3235 1266 3269
rect 1232 3163 1266 3197
rect 1232 3091 1266 3125
rect 1232 3019 1266 3053
rect 1232 2947 1266 2981
rect 1232 2875 1266 2909
rect 1232 2803 1266 2837
rect 1232 2731 1266 2765
rect 1232 2659 1266 2693
rect 1232 2587 1266 2621
rect 1232 2515 1266 2549
rect 1232 2443 1266 2477
rect 1232 2371 1266 2405
rect 1232 2299 1266 2333
rect 1232 2227 1266 2261
rect 1232 2155 1266 2189
rect 1232 2083 1266 2117
rect 1232 2011 1266 2045
rect 1232 1939 1266 1973
rect 1232 1867 1266 1901
rect 1232 1795 1266 1829
rect 1232 1723 1266 1757
rect 1232 1651 1266 1685
rect 1232 1579 1266 1613
rect 1232 1507 1266 1541
rect 1232 1435 1266 1469
rect 1232 1363 1266 1397
rect 1232 1291 1266 1325
rect 1232 1219 1266 1253
rect 1232 1147 1266 1181
rect 1232 1075 1266 1109
rect 1232 1003 1266 1037
rect 1232 931 1266 965
rect 1232 859 1266 893
rect 1232 787 1266 821
rect 1232 715 1266 749
rect 1232 643 1266 677
rect 1232 571 1266 605
rect 1232 499 1266 533
rect 1232 427 1266 461
rect 1232 355 1266 389
rect 1232 283 1266 317
rect 1232 211 1266 245
rect 1232 139 1266 173
rect 1232 67 1266 101
rect -1116 -77 -1082 -43
rect -1116 -149 -1082 -115
rect -1116 -221 -1082 -187
rect -1116 -293 -1082 -259
rect -1116 -365 -1082 -331
rect -1116 -437 -1082 -403
rect -1116 -509 -1082 -475
rect -1116 -581 -1082 -547
rect -1116 -653 -1082 -619
rect 1232 -5 1266 29
rect 1232 -77 1266 -43
rect 1232 -149 1266 -115
rect 1232 -221 1266 -187
rect 1232 -293 1266 -259
rect 1232 -365 1266 -331
rect 1232 -437 1266 -403
rect 1232 -509 1266 -475
rect 1232 -581 1266 -547
rect -1116 -725 -1082 -691
rect -1116 -797 -1082 -763
rect -1116 -869 -1082 -835
rect -280 -693 -246 -659
rect -206 -693 -172 -659
rect -132 -693 -98 -659
rect -58 -693 -24 -659
rect 16 -693 50 -659
rect 90 -693 124 -659
rect 164 -693 198 -659
rect 238 -693 272 -659
rect 312 -693 346 -659
rect 386 -693 420 -659
rect -280 -767 -246 -733
rect -206 -767 -172 -733
rect -132 -767 -98 -733
rect -58 -767 -24 -733
rect 16 -767 50 -733
rect 90 -767 124 -733
rect 164 -767 198 -733
rect 238 -767 272 -733
rect 312 -767 346 -733
rect 386 -767 420 -733
rect -280 -841 -246 -807
rect -206 -841 -172 -807
rect -132 -841 -98 -807
rect -58 -841 -24 -807
rect 16 -841 50 -807
rect 90 -841 124 -807
rect 164 -841 198 -807
rect 238 -841 272 -807
rect 312 -841 346 -807
rect 386 -841 420 -807
rect 1232 -653 1266 -619
rect 1232 -725 1266 -691
rect 1232 -797 1266 -763
rect -1116 -941 -1082 -907
rect -1116 -1013 -1082 -979
rect -1116 -1085 -1082 -1051
rect 1232 -869 1266 -835
rect 1232 -941 1266 -907
rect 1232 -1013 1266 -979
rect 1232 -1085 1266 -1051
rect -988 -1158 -954 -1124
rect -916 -1158 -882 -1124
rect -844 -1158 -810 -1124
rect -772 -1158 -738 -1124
rect -700 -1158 -666 -1124
rect -628 -1158 -594 -1124
rect -556 -1158 -522 -1124
rect -484 -1158 -450 -1124
rect -412 -1158 -378 -1124
rect -340 -1158 -306 -1124
rect -268 -1158 -234 -1124
rect -196 -1158 -162 -1124
rect -124 -1158 -90 -1124
rect -52 -1158 -18 -1124
rect 20 -1158 54 -1124
rect 92 -1158 126 -1124
rect 164 -1158 198 -1124
rect 236 -1158 270 -1124
rect 308 -1158 342 -1124
rect 380 -1158 414 -1124
rect 452 -1158 486 -1124
rect 524 -1158 558 -1124
rect 596 -1158 630 -1124
rect 668 -1158 702 -1124
rect 740 -1158 774 -1124
rect 812 -1158 846 -1124
rect 884 -1158 918 -1124
rect 956 -1158 990 -1124
rect 1028 -1158 1062 -1124
rect 1100 -1158 1134 -1124
<< metal1 >>
rect -1140 7158 1290 7182
rect -1140 7124 -988 7158
rect -954 7124 -916 7158
rect -882 7124 -844 7158
rect -810 7124 -772 7158
rect -738 7124 -700 7158
rect -666 7124 -628 7158
rect -594 7124 -556 7158
rect -522 7124 -484 7158
rect -450 7124 -412 7158
rect -378 7124 -340 7158
rect -306 7124 -268 7158
rect -234 7124 -196 7158
rect -162 7124 -124 7158
rect -90 7124 -52 7158
rect -18 7124 20 7158
rect 54 7124 92 7158
rect 126 7124 164 7158
rect 198 7124 236 7158
rect 270 7124 308 7158
rect 342 7124 380 7158
rect 414 7124 452 7158
rect 486 7124 524 7158
rect 558 7124 596 7158
rect 630 7124 668 7158
rect 702 7124 740 7158
rect 774 7124 812 7158
rect 846 7124 884 7158
rect 918 7124 956 7158
rect 990 7124 1028 7158
rect 1062 7124 1100 7158
rect 1134 7124 1290 7158
rect -1140 7100 1290 7124
rect -1140 7085 -1058 7100
rect -1140 7051 -1116 7085
rect -1082 7051 -1058 7085
rect -1140 7013 -1058 7051
rect -1140 6979 -1116 7013
rect -1082 6979 -1058 7013
rect -1140 6941 -1058 6979
rect -1140 6907 -1116 6941
rect -1082 6907 -1058 6941
rect -1140 6869 -1058 6907
rect -1140 6835 -1116 6869
rect -1082 6835 -1058 6869
rect -1140 6797 -1058 6835
rect -1140 6763 -1116 6797
rect -1082 6763 -1058 6797
rect -1140 6725 -1058 6763
rect -1140 6691 -1116 6725
rect -1082 6691 -1058 6725
rect -1140 6653 -1058 6691
rect -1140 6619 -1116 6653
rect -1082 6619 -1058 6653
rect -1140 6581 -1058 6619
rect -1140 6547 -1116 6581
rect -1082 6547 -1058 6581
rect -1140 6509 -1058 6547
rect -1140 6475 -1116 6509
rect -1082 6475 -1058 6509
rect -1140 6437 -1058 6475
rect -1140 6403 -1116 6437
rect -1082 6403 -1058 6437
rect -1140 6365 -1058 6403
rect -1140 6331 -1116 6365
rect -1082 6331 -1058 6365
rect -1140 6293 -1058 6331
rect -1140 6259 -1116 6293
rect -1082 6259 -1058 6293
rect -1140 6221 -1058 6259
rect -1140 6187 -1116 6221
rect -1082 6187 -1058 6221
rect -1140 6149 -1058 6187
rect -1140 6115 -1116 6149
rect -1082 6115 -1058 6149
rect -1140 6077 -1058 6115
rect -1140 6043 -1116 6077
rect -1082 6043 -1058 6077
rect -1140 6005 -1058 6043
rect -1140 5971 -1116 6005
rect -1082 5971 -1058 6005
rect 1208 7085 1290 7100
rect 1208 7051 1232 7085
rect 1266 7051 1290 7085
rect 1208 7013 1290 7051
rect 1208 6979 1232 7013
rect 1266 6979 1290 7013
rect 1208 6941 1290 6979
rect 1208 6907 1232 6941
rect 1266 6907 1290 6941
rect 1208 6869 1290 6907
rect 1208 6835 1232 6869
rect 1266 6835 1290 6869
rect 1208 6797 1290 6835
rect 1208 6763 1232 6797
rect 1266 6763 1290 6797
rect 1208 6725 1290 6763
rect 1208 6691 1232 6725
rect 1266 6691 1290 6725
rect 1208 6653 1290 6691
rect 1208 6619 1232 6653
rect 1266 6619 1290 6653
rect 1208 6581 1290 6619
rect 1208 6547 1232 6581
rect 1266 6547 1290 6581
rect 1208 6509 1290 6547
rect 1208 6475 1232 6509
rect 1266 6475 1290 6509
rect 1208 6437 1290 6475
rect 1208 6403 1232 6437
rect 1266 6403 1290 6437
rect 1208 6365 1290 6403
rect 1208 6331 1232 6365
rect 1266 6331 1290 6365
rect 1208 6293 1290 6331
rect 1208 6259 1232 6293
rect 1266 6259 1290 6293
rect 1208 6221 1290 6259
rect 1208 6187 1232 6221
rect 1266 6187 1290 6221
rect 1208 6149 1290 6187
rect 1208 6115 1232 6149
rect 1266 6115 1290 6149
rect 1208 6077 1290 6115
rect 1208 6043 1232 6077
rect 1266 6043 1290 6077
rect 1208 6005 1290 6043
rect -1140 5933 -1058 5971
rect -1140 5899 -1116 5933
rect -1082 5899 -1058 5933
rect -1140 5861 -1058 5899
rect -1140 5827 -1116 5861
rect -1082 5827 -1058 5861
rect -1140 5789 -1058 5827
rect -1140 5755 -1116 5789
rect -1082 5755 -1058 5789
rect -1140 5717 -1058 5755
rect -1140 5683 -1116 5717
rect -1082 5683 -1058 5717
rect -1140 5645 -1058 5683
rect -1140 5611 -1116 5645
rect -1082 5611 -1058 5645
rect -1140 5573 -1058 5611
rect -1140 5539 -1116 5573
rect -1082 5539 -1058 5573
rect -1140 5501 -1058 5539
rect -1140 5467 -1116 5501
rect -1082 5467 -1058 5501
rect -1140 5429 -1058 5467
rect -1140 5395 -1116 5429
rect -1082 5395 -1058 5429
rect -1140 5357 -1058 5395
rect -1140 5323 -1116 5357
rect -1082 5323 -1058 5357
rect -1140 5285 -1058 5323
rect -1140 5251 -1116 5285
rect -1082 5251 -1058 5285
rect -1140 5213 -1058 5251
rect -1140 5179 -1116 5213
rect -1082 5179 -1058 5213
rect -1140 5141 -1058 5179
rect -1140 5107 -1116 5141
rect -1082 5107 -1058 5141
rect -1140 5069 -1058 5107
rect -1140 5035 -1116 5069
rect -1082 5035 -1058 5069
rect -1140 4997 -1058 5035
rect -1140 4963 -1116 4997
rect -1082 4963 -1058 4997
rect -1140 4925 -1058 4963
rect -1140 4891 -1116 4925
rect -1082 4891 -1058 4925
rect -1140 4853 -1058 4891
rect -1140 4819 -1116 4853
rect -1082 4819 -1058 4853
rect -1140 4781 -1058 4819
rect -1140 4747 -1116 4781
rect -1082 4747 -1058 4781
rect -1140 4709 -1058 4747
rect -1140 4675 -1116 4709
rect -1082 4675 -1058 4709
rect -1140 4637 -1058 4675
rect -1140 4603 -1116 4637
rect -1082 4603 -1058 4637
rect -1140 4565 -1058 4603
rect -1140 4531 -1116 4565
rect -1082 4531 -1058 4565
rect -1140 4493 -1058 4531
rect -1140 4459 -1116 4493
rect -1082 4459 -1058 4493
rect -1140 4421 -1058 4459
rect -1140 4387 -1116 4421
rect -1082 4387 -1058 4421
rect -1140 4349 -1058 4387
rect -1140 4315 -1116 4349
rect -1082 4315 -1058 4349
rect -1140 4277 -1058 4315
rect -1140 4243 -1116 4277
rect -1082 4243 -1058 4277
rect -1140 4205 -1058 4243
rect -1140 4171 -1116 4205
rect -1082 4171 -1058 4205
rect -1140 4133 -1058 4171
rect -1140 4099 -1116 4133
rect -1082 4099 -1058 4133
rect -1140 4061 -1058 4099
rect -1140 4027 -1116 4061
rect -1082 4027 -1058 4061
rect -1140 3989 -1058 4027
rect -1140 3955 -1116 3989
rect -1082 3955 -1058 3989
rect -1140 3917 -1058 3955
rect -1140 3883 -1116 3917
rect -1082 3883 -1058 3917
rect -1140 3845 -1058 3883
rect -1140 3811 -1116 3845
rect -1082 3811 -1058 3845
rect -1140 3773 -1058 3811
rect -1140 3739 -1116 3773
rect -1082 3739 -1058 3773
rect -1140 3701 -1058 3739
rect -1140 3667 -1116 3701
rect -1082 3667 -1058 3701
rect -1140 3629 -1058 3667
rect -1140 3595 -1116 3629
rect -1082 3595 -1058 3629
rect -1140 3557 -1058 3595
rect -1140 3523 -1116 3557
rect -1082 3523 -1058 3557
rect -1140 3485 -1058 3523
rect -1140 3451 -1116 3485
rect -1082 3451 -1058 3485
rect -1140 3413 -1058 3451
rect -1140 3379 -1116 3413
rect -1082 3379 -1058 3413
rect -1140 3341 -1058 3379
rect -1140 3307 -1116 3341
rect -1082 3307 -1058 3341
rect -1140 3269 -1058 3307
rect -1140 3235 -1116 3269
rect -1082 3235 -1058 3269
rect -1140 3197 -1058 3235
rect -1140 3163 -1116 3197
rect -1082 3163 -1058 3197
rect -1140 3125 -1058 3163
rect -1140 3091 -1116 3125
rect -1082 3091 -1058 3125
rect -1140 3053 -1058 3091
rect -1140 3019 -1116 3053
rect -1082 3019 -1058 3053
rect -1140 2981 -1058 3019
rect -1140 2947 -1116 2981
rect -1082 2947 -1058 2981
rect -1140 2909 -1058 2947
rect -1140 2875 -1116 2909
rect -1082 2875 -1058 2909
rect -1140 2837 -1058 2875
rect -1140 2803 -1116 2837
rect -1082 2803 -1058 2837
rect -1140 2765 -1058 2803
rect -1140 2731 -1116 2765
rect -1082 2731 -1058 2765
rect -1140 2693 -1058 2731
rect -1140 2659 -1116 2693
rect -1082 2659 -1058 2693
rect -1140 2621 -1058 2659
rect -1140 2587 -1116 2621
rect -1082 2587 -1058 2621
rect -1140 2549 -1058 2587
rect -1140 2515 -1116 2549
rect -1082 2515 -1058 2549
rect -1140 2477 -1058 2515
rect -1140 2443 -1116 2477
rect -1082 2443 -1058 2477
rect -1140 2405 -1058 2443
rect -1140 2371 -1116 2405
rect -1082 2371 -1058 2405
rect -1140 2333 -1058 2371
rect -1140 2299 -1116 2333
rect -1082 2299 -1058 2333
rect -1140 2261 -1058 2299
rect -1140 2227 -1116 2261
rect -1082 2227 -1058 2261
rect -1140 2189 -1058 2227
rect -1140 2155 -1116 2189
rect -1082 2155 -1058 2189
rect -1140 2117 -1058 2155
rect -1140 2083 -1116 2117
rect -1082 2083 -1058 2117
rect -1140 2045 -1058 2083
rect -1140 2011 -1116 2045
rect -1082 2011 -1058 2045
rect -1140 1973 -1058 2011
rect -1140 1939 -1116 1973
rect -1082 1939 -1058 1973
rect -1140 1901 -1058 1939
rect -1140 1867 -1116 1901
rect -1082 1867 -1058 1901
rect -1140 1829 -1058 1867
rect -1140 1795 -1116 1829
rect -1082 1795 -1058 1829
rect -1140 1757 -1058 1795
rect -1140 1723 -1116 1757
rect -1082 1723 -1058 1757
rect -1140 1685 -1058 1723
rect -1140 1651 -1116 1685
rect -1082 1651 -1058 1685
rect -1140 1613 -1058 1651
rect -1140 1579 -1116 1613
rect -1082 1579 -1058 1613
rect -1140 1541 -1058 1579
rect -1140 1507 -1116 1541
rect -1082 1507 -1058 1541
rect -1140 1469 -1058 1507
rect -1140 1435 -1116 1469
rect -1082 1435 -1058 1469
rect -1140 1397 -1058 1435
rect -1140 1363 -1116 1397
rect -1082 1363 -1058 1397
rect -1140 1325 -1058 1363
rect -1140 1291 -1116 1325
rect -1082 1291 -1058 1325
rect -1140 1253 -1058 1291
rect -1140 1219 -1116 1253
rect -1082 1219 -1058 1253
rect -1140 1181 -1058 1219
rect -1140 1147 -1116 1181
rect -1082 1147 -1058 1181
rect -1140 1109 -1058 1147
rect -1140 1075 -1116 1109
rect -1082 1075 -1058 1109
rect -1140 1037 -1058 1075
rect -1140 1003 -1116 1037
rect -1082 1003 -1058 1037
rect -1140 965 -1058 1003
rect -1140 931 -1116 965
rect -1082 931 -1058 965
rect -1140 893 -1058 931
rect -1140 859 -1116 893
rect -1082 859 -1058 893
rect -1140 821 -1058 859
rect -1140 787 -1116 821
rect -1082 787 -1058 821
rect -1140 749 -1058 787
rect -1140 715 -1116 749
rect -1082 715 -1058 749
rect -1140 677 -1058 715
rect -1140 643 -1116 677
rect -1082 643 -1058 677
rect -1140 605 -1058 643
rect -1140 571 -1116 605
rect -1082 571 -1058 605
rect -1140 533 -1058 571
rect -1140 499 -1116 533
rect -1082 499 -1058 533
rect -1140 461 -1058 499
rect -1140 427 -1116 461
rect -1082 427 -1058 461
rect -1140 389 -1058 427
rect -1140 355 -1116 389
rect -1082 355 -1058 389
rect -1140 317 -1058 355
rect -1140 283 -1116 317
rect -1082 283 -1058 317
rect -1140 245 -1058 283
rect -1140 211 -1116 245
rect -1082 211 -1058 245
rect -1140 173 -1058 211
rect -1140 139 -1116 173
rect -1082 139 -1058 173
rect -1140 101 -1058 139
rect -1140 67 -1116 101
rect -1082 67 -1058 101
rect -1140 29 -1058 67
rect -1140 -5 -1116 29
rect -1082 -5 -1058 29
rect -958 5969 -900 5981
rect -958 5935 -946 5969
rect -912 5935 -900 5969
rect 1050 5969 1108 5981
rect -958 5897 -900 5935
rect -958 5863 -946 5897
rect -912 5863 -900 5897
rect -958 5825 -900 5863
rect -958 5791 -946 5825
rect -912 5791 -900 5825
rect -958 5753 -900 5791
rect -958 5719 -946 5753
rect -912 5719 -900 5753
rect -958 5681 -900 5719
rect -958 5647 -946 5681
rect -912 5647 -900 5681
rect -958 5609 -900 5647
rect -958 5575 -946 5609
rect -912 5575 -900 5609
rect -958 5537 -900 5575
rect -958 5503 -946 5537
rect -912 5503 -900 5537
rect -958 5465 -900 5503
rect -958 5431 -946 5465
rect -912 5431 -900 5465
rect -958 5393 -900 5431
rect -958 5359 -946 5393
rect -912 5359 -900 5393
rect -958 5321 -900 5359
rect -958 5287 -946 5321
rect -912 5287 -900 5321
rect -958 5249 -900 5287
rect -958 5215 -946 5249
rect -912 5215 -900 5249
rect -958 5177 -900 5215
rect -958 5143 -946 5177
rect -912 5143 -900 5177
rect -958 5105 -900 5143
rect -958 5071 -946 5105
rect -912 5071 -900 5105
rect -958 5033 -900 5071
rect -958 4999 -946 5033
rect -912 4999 -900 5033
rect -958 4961 -900 4999
rect -958 4927 -946 4961
rect -912 4927 -900 4961
rect -958 4889 -900 4927
rect -958 4855 -946 4889
rect -912 4855 -900 4889
rect -958 4817 -900 4855
rect -958 4783 -946 4817
rect -912 4783 -900 4817
rect -958 4745 -900 4783
rect -958 4711 -946 4745
rect -912 4711 -900 4745
rect -958 4673 -900 4711
rect -958 4639 -946 4673
rect -912 4639 -900 4673
rect -958 4601 -900 4639
rect -958 4567 -946 4601
rect -912 4567 -900 4601
rect -958 4529 -900 4567
rect -958 4495 -946 4529
rect -912 4495 -900 4529
rect -958 4457 -900 4495
rect -958 4423 -946 4457
rect -912 4423 -900 4457
rect -958 4385 -900 4423
rect -958 4351 -946 4385
rect -912 4351 -900 4385
rect -958 4313 -900 4351
rect -958 4279 -946 4313
rect -912 4279 -900 4313
rect -958 4241 -900 4279
rect -958 4207 -946 4241
rect -912 4207 -900 4241
rect -958 4169 -900 4207
rect -958 4135 -946 4169
rect -912 4135 -900 4169
rect -958 4097 -900 4135
rect -958 4063 -946 4097
rect -912 4063 -900 4097
rect -958 4025 -900 4063
rect -958 3991 -946 4025
rect -912 3991 -900 4025
rect -958 3953 -900 3991
rect -958 3919 -946 3953
rect -912 3919 -900 3953
rect -958 3881 -900 3919
rect -958 3847 -946 3881
rect -912 3847 -900 3881
rect -958 3809 -900 3847
rect -958 3775 -946 3809
rect -912 3775 -900 3809
rect -958 3737 -900 3775
rect -958 3703 -946 3737
rect -912 3703 -900 3737
rect -958 3665 -900 3703
rect -958 3631 -946 3665
rect -912 3631 -900 3665
rect -958 3593 -900 3631
rect -958 3559 -946 3593
rect -912 3559 -900 3593
rect -958 3521 -900 3559
rect -958 3487 -946 3521
rect -912 3487 -900 3521
rect -958 3449 -900 3487
rect -958 3415 -946 3449
rect -912 3415 -900 3449
rect -958 3377 -900 3415
rect -958 3343 -946 3377
rect -912 3343 -900 3377
rect -958 3305 -900 3343
rect -958 3271 -946 3305
rect -912 3271 -900 3305
rect -958 3233 -900 3271
rect -958 3199 -946 3233
rect -912 3199 -900 3233
rect -958 3161 -900 3199
rect -958 3127 -946 3161
rect -912 3127 -900 3161
rect -958 3089 -900 3127
rect -958 3055 -946 3089
rect -912 3055 -900 3089
rect -958 3017 -900 3055
rect -958 2983 -946 3017
rect -912 2983 -900 3017
rect -958 2945 -900 2983
rect -958 2911 -946 2945
rect -912 2911 -900 2945
rect -958 2873 -900 2911
rect -958 2839 -946 2873
rect -912 2839 -900 2873
rect -958 2801 -900 2839
rect -958 2767 -946 2801
rect -912 2767 -900 2801
rect -958 2729 -900 2767
rect -958 2695 -946 2729
rect -912 2695 -900 2729
rect -958 2657 -900 2695
rect -958 2623 -946 2657
rect -912 2623 -900 2657
rect -958 2585 -900 2623
rect -958 2551 -946 2585
rect -912 2551 -900 2585
rect -958 2513 -900 2551
rect -958 2479 -946 2513
rect -912 2479 -900 2513
rect -958 2441 -900 2479
rect -958 2407 -946 2441
rect -912 2407 -900 2441
rect -958 2369 -900 2407
rect -958 2335 -946 2369
rect -912 2335 -900 2369
rect -958 2297 -900 2335
rect -958 2263 -946 2297
rect -912 2263 -900 2297
rect -958 2225 -900 2263
rect -958 2191 -946 2225
rect -912 2191 -900 2225
rect -958 2153 -900 2191
rect -958 2119 -946 2153
rect -912 2119 -900 2153
rect -958 2081 -900 2119
rect -958 2047 -946 2081
rect -912 2047 -900 2081
rect -958 2009 -900 2047
rect -958 1975 -946 2009
rect -912 1975 -900 2009
rect -958 1937 -900 1975
rect -958 1903 -946 1937
rect -912 1903 -900 1937
rect -958 1865 -900 1903
rect -958 1831 -946 1865
rect -912 1831 -900 1865
rect -958 1793 -900 1831
rect -958 1759 -946 1793
rect -912 1759 -900 1793
rect -958 1721 -900 1759
rect -958 1687 -946 1721
rect -912 1687 -900 1721
rect -958 1649 -900 1687
rect -958 1615 -946 1649
rect -912 1615 -900 1649
rect -958 1577 -900 1615
rect -958 1543 -946 1577
rect -912 1543 -900 1577
rect -958 1505 -900 1543
rect -958 1471 -946 1505
rect -912 1471 -900 1505
rect -958 1433 -900 1471
rect -958 1399 -946 1433
rect -912 1399 -900 1433
rect -958 1361 -900 1399
rect -958 1327 -946 1361
rect -912 1327 -900 1361
rect -958 1289 -900 1327
rect -958 1255 -946 1289
rect -912 1255 -900 1289
rect -958 1217 -900 1255
rect -958 1183 -946 1217
rect -912 1183 -900 1217
rect -958 1145 -900 1183
rect -958 1111 -946 1145
rect -912 1111 -900 1145
rect -958 1073 -900 1111
rect -958 1039 -946 1073
rect -912 1039 -900 1073
rect -958 1001 -900 1039
rect -958 967 -946 1001
rect -912 967 -900 1001
rect -958 929 -900 967
rect -958 895 -946 929
rect -912 895 -900 929
rect -958 857 -900 895
rect -958 823 -946 857
rect -912 823 -900 857
rect -958 785 -900 823
rect -958 751 -946 785
rect -912 751 -900 785
rect -958 713 -900 751
rect -958 679 -946 713
rect -912 679 -900 713
rect -958 641 -900 679
rect -958 607 -946 641
rect -912 607 -900 641
rect -958 569 -900 607
rect -958 535 -946 569
rect -912 535 -900 569
rect -958 497 -900 535
rect -958 463 -946 497
rect -912 463 -900 497
rect -958 425 -900 463
rect -958 391 -946 425
rect -912 391 -900 425
rect -958 353 -900 391
rect -958 319 -946 353
rect -912 319 -900 353
rect -958 281 -900 319
rect -958 247 -946 281
rect -912 247 -900 281
rect -958 209 -900 247
rect -958 175 -946 209
rect -912 175 -900 209
rect -958 137 -900 175
rect -958 103 -946 137
rect -912 103 -900 137
rect -958 65 -900 103
rect -958 31 -946 65
rect -912 31 -900 65
rect 10 5939 140 5945
rect 10 63 17 5939
rect 133 63 140 5939
rect 10 55 140 63
rect 1050 5935 1062 5969
rect 1096 5935 1108 5969
rect 1050 5897 1108 5935
rect 1050 5863 1062 5897
rect 1096 5863 1108 5897
rect 1050 5825 1108 5863
rect 1050 5791 1062 5825
rect 1096 5791 1108 5825
rect 1050 5753 1108 5791
rect 1050 5719 1062 5753
rect 1096 5719 1108 5753
rect 1050 5681 1108 5719
rect 1050 5647 1062 5681
rect 1096 5647 1108 5681
rect 1050 5609 1108 5647
rect 1050 5575 1062 5609
rect 1096 5575 1108 5609
rect 1050 5537 1108 5575
rect 1050 5503 1062 5537
rect 1096 5503 1108 5537
rect 1050 5465 1108 5503
rect 1050 5431 1062 5465
rect 1096 5431 1108 5465
rect 1050 5393 1108 5431
rect 1050 5359 1062 5393
rect 1096 5359 1108 5393
rect 1050 5321 1108 5359
rect 1050 5287 1062 5321
rect 1096 5287 1108 5321
rect 1050 5249 1108 5287
rect 1050 5215 1062 5249
rect 1096 5215 1108 5249
rect 1050 5177 1108 5215
rect 1050 5143 1062 5177
rect 1096 5143 1108 5177
rect 1050 5105 1108 5143
rect 1050 5071 1062 5105
rect 1096 5071 1108 5105
rect 1050 5033 1108 5071
rect 1050 4999 1062 5033
rect 1096 4999 1108 5033
rect 1050 4961 1108 4999
rect 1050 4927 1062 4961
rect 1096 4927 1108 4961
rect 1050 4889 1108 4927
rect 1050 4855 1062 4889
rect 1096 4855 1108 4889
rect 1050 4817 1108 4855
rect 1050 4783 1062 4817
rect 1096 4783 1108 4817
rect 1050 4745 1108 4783
rect 1050 4711 1062 4745
rect 1096 4711 1108 4745
rect 1050 4673 1108 4711
rect 1050 4639 1062 4673
rect 1096 4639 1108 4673
rect 1050 4601 1108 4639
rect 1050 4567 1062 4601
rect 1096 4567 1108 4601
rect 1050 4529 1108 4567
rect 1050 4495 1062 4529
rect 1096 4495 1108 4529
rect 1050 4457 1108 4495
rect 1050 4423 1062 4457
rect 1096 4423 1108 4457
rect 1050 4385 1108 4423
rect 1050 4351 1062 4385
rect 1096 4351 1108 4385
rect 1050 4313 1108 4351
rect 1050 4279 1062 4313
rect 1096 4279 1108 4313
rect 1050 4241 1108 4279
rect 1050 4207 1062 4241
rect 1096 4207 1108 4241
rect 1050 4169 1108 4207
rect 1050 4135 1062 4169
rect 1096 4135 1108 4169
rect 1050 4097 1108 4135
rect 1050 4063 1062 4097
rect 1096 4063 1108 4097
rect 1050 4025 1108 4063
rect 1050 3991 1062 4025
rect 1096 3991 1108 4025
rect 1050 3953 1108 3991
rect 1050 3919 1062 3953
rect 1096 3919 1108 3953
rect 1050 3881 1108 3919
rect 1050 3847 1062 3881
rect 1096 3847 1108 3881
rect 1050 3809 1108 3847
rect 1050 3775 1062 3809
rect 1096 3775 1108 3809
rect 1050 3737 1108 3775
rect 1050 3703 1062 3737
rect 1096 3703 1108 3737
rect 1050 3665 1108 3703
rect 1050 3631 1062 3665
rect 1096 3631 1108 3665
rect 1050 3593 1108 3631
rect 1050 3559 1062 3593
rect 1096 3559 1108 3593
rect 1050 3521 1108 3559
rect 1050 3487 1062 3521
rect 1096 3487 1108 3521
rect 1050 3449 1108 3487
rect 1050 3415 1062 3449
rect 1096 3415 1108 3449
rect 1050 3377 1108 3415
rect 1050 3343 1062 3377
rect 1096 3343 1108 3377
rect 1050 3305 1108 3343
rect 1050 3271 1062 3305
rect 1096 3271 1108 3305
rect 1050 3233 1108 3271
rect 1050 3199 1062 3233
rect 1096 3199 1108 3233
rect 1050 3161 1108 3199
rect 1050 3127 1062 3161
rect 1096 3127 1108 3161
rect 1050 3089 1108 3127
rect 1050 3055 1062 3089
rect 1096 3055 1108 3089
rect 1050 3017 1108 3055
rect 1050 2983 1062 3017
rect 1096 2983 1108 3017
rect 1050 2945 1108 2983
rect 1050 2911 1062 2945
rect 1096 2911 1108 2945
rect 1050 2873 1108 2911
rect 1050 2839 1062 2873
rect 1096 2839 1108 2873
rect 1050 2801 1108 2839
rect 1050 2767 1062 2801
rect 1096 2767 1108 2801
rect 1050 2729 1108 2767
rect 1050 2695 1062 2729
rect 1096 2695 1108 2729
rect 1050 2657 1108 2695
rect 1050 2623 1062 2657
rect 1096 2623 1108 2657
rect 1050 2585 1108 2623
rect 1050 2551 1062 2585
rect 1096 2551 1108 2585
rect 1050 2513 1108 2551
rect 1050 2479 1062 2513
rect 1096 2479 1108 2513
rect 1050 2441 1108 2479
rect 1050 2407 1062 2441
rect 1096 2407 1108 2441
rect 1050 2369 1108 2407
rect 1050 2335 1062 2369
rect 1096 2335 1108 2369
rect 1050 2297 1108 2335
rect 1050 2263 1062 2297
rect 1096 2263 1108 2297
rect 1050 2225 1108 2263
rect 1050 2191 1062 2225
rect 1096 2191 1108 2225
rect 1050 2153 1108 2191
rect 1050 2119 1062 2153
rect 1096 2119 1108 2153
rect 1050 2081 1108 2119
rect 1050 2047 1062 2081
rect 1096 2047 1108 2081
rect 1050 2009 1108 2047
rect 1050 1975 1062 2009
rect 1096 1975 1108 2009
rect 1050 1937 1108 1975
rect 1050 1903 1062 1937
rect 1096 1903 1108 1937
rect 1050 1865 1108 1903
rect 1050 1831 1062 1865
rect 1096 1831 1108 1865
rect 1050 1793 1108 1831
rect 1050 1759 1062 1793
rect 1096 1759 1108 1793
rect 1050 1721 1108 1759
rect 1050 1687 1062 1721
rect 1096 1687 1108 1721
rect 1050 1649 1108 1687
rect 1050 1615 1062 1649
rect 1096 1615 1108 1649
rect 1050 1577 1108 1615
rect 1050 1543 1062 1577
rect 1096 1543 1108 1577
rect 1050 1505 1108 1543
rect 1050 1471 1062 1505
rect 1096 1471 1108 1505
rect 1050 1433 1108 1471
rect 1050 1399 1062 1433
rect 1096 1399 1108 1433
rect 1050 1361 1108 1399
rect 1050 1327 1062 1361
rect 1096 1327 1108 1361
rect 1050 1289 1108 1327
rect 1050 1255 1062 1289
rect 1096 1255 1108 1289
rect 1050 1217 1108 1255
rect 1050 1183 1062 1217
rect 1096 1183 1108 1217
rect 1050 1145 1108 1183
rect 1050 1111 1062 1145
rect 1096 1111 1108 1145
rect 1050 1073 1108 1111
rect 1050 1039 1062 1073
rect 1096 1039 1108 1073
rect 1050 1001 1108 1039
rect 1050 967 1062 1001
rect 1096 967 1108 1001
rect 1050 929 1108 967
rect 1050 895 1062 929
rect 1096 895 1108 929
rect 1050 857 1108 895
rect 1050 823 1062 857
rect 1096 823 1108 857
rect 1050 785 1108 823
rect 1050 751 1062 785
rect 1096 751 1108 785
rect 1050 713 1108 751
rect 1050 679 1062 713
rect 1096 679 1108 713
rect 1050 641 1108 679
rect 1050 607 1062 641
rect 1096 607 1108 641
rect 1050 569 1108 607
rect 1050 535 1062 569
rect 1096 535 1108 569
rect 1050 497 1108 535
rect 1050 463 1062 497
rect 1096 463 1108 497
rect 1050 425 1108 463
rect 1050 391 1062 425
rect 1096 391 1108 425
rect 1050 353 1108 391
rect 1050 319 1062 353
rect 1096 319 1108 353
rect 1050 281 1108 319
rect 1050 247 1062 281
rect 1096 247 1108 281
rect 1050 209 1108 247
rect 1050 175 1062 209
rect 1096 175 1108 209
rect 1050 137 1108 175
rect 1050 103 1062 137
rect 1096 103 1108 137
rect 1050 65 1108 103
rect -958 19 -900 31
rect 1050 31 1062 65
rect 1096 31 1108 65
rect 1050 19 1108 31
rect 1208 5971 1232 6005
rect 1266 5971 1290 6005
rect 1208 5933 1290 5971
rect 1208 5899 1232 5933
rect 1266 5899 1290 5933
rect 1208 5861 1290 5899
rect 1208 5827 1232 5861
rect 1266 5827 1290 5861
rect 1208 5789 1290 5827
rect 1208 5755 1232 5789
rect 1266 5755 1290 5789
rect 1208 5717 1290 5755
rect 1208 5683 1232 5717
rect 1266 5683 1290 5717
rect 1208 5645 1290 5683
rect 1208 5611 1232 5645
rect 1266 5611 1290 5645
rect 1208 5573 1290 5611
rect 1208 5539 1232 5573
rect 1266 5539 1290 5573
rect 1208 5501 1290 5539
rect 1208 5467 1232 5501
rect 1266 5467 1290 5501
rect 1208 5429 1290 5467
rect 1208 5395 1232 5429
rect 1266 5395 1290 5429
rect 1208 5357 1290 5395
rect 1208 5323 1232 5357
rect 1266 5323 1290 5357
rect 1208 5285 1290 5323
rect 1208 5251 1232 5285
rect 1266 5251 1290 5285
rect 1208 5213 1290 5251
rect 1208 5179 1232 5213
rect 1266 5179 1290 5213
rect 1208 5141 1290 5179
rect 1208 5107 1232 5141
rect 1266 5107 1290 5141
rect 1208 5069 1290 5107
rect 1208 5035 1232 5069
rect 1266 5035 1290 5069
rect 1208 4997 1290 5035
rect 1208 4963 1232 4997
rect 1266 4963 1290 4997
rect 1208 4925 1290 4963
rect 1208 4891 1232 4925
rect 1266 4891 1290 4925
rect 1208 4853 1290 4891
rect 1208 4819 1232 4853
rect 1266 4819 1290 4853
rect 1208 4781 1290 4819
rect 1208 4747 1232 4781
rect 1266 4747 1290 4781
rect 1208 4709 1290 4747
rect 1208 4675 1232 4709
rect 1266 4675 1290 4709
rect 1208 4637 1290 4675
rect 1208 4603 1232 4637
rect 1266 4603 1290 4637
rect 1208 4565 1290 4603
rect 1208 4531 1232 4565
rect 1266 4531 1290 4565
rect 1208 4493 1290 4531
rect 1208 4459 1232 4493
rect 1266 4459 1290 4493
rect 1208 4421 1290 4459
rect 1208 4387 1232 4421
rect 1266 4387 1290 4421
rect 1208 4349 1290 4387
rect 1208 4315 1232 4349
rect 1266 4315 1290 4349
rect 1208 4277 1290 4315
rect 1208 4243 1232 4277
rect 1266 4243 1290 4277
rect 1208 4205 1290 4243
rect 1208 4171 1232 4205
rect 1266 4171 1290 4205
rect 1208 4133 1290 4171
rect 1208 4099 1232 4133
rect 1266 4099 1290 4133
rect 1208 4061 1290 4099
rect 1208 4027 1232 4061
rect 1266 4027 1290 4061
rect 1208 3989 1290 4027
rect 1208 3955 1232 3989
rect 1266 3955 1290 3989
rect 1208 3917 1290 3955
rect 1208 3883 1232 3917
rect 1266 3883 1290 3917
rect 1208 3845 1290 3883
rect 1208 3811 1232 3845
rect 1266 3811 1290 3845
rect 1208 3773 1290 3811
rect 1208 3739 1232 3773
rect 1266 3739 1290 3773
rect 1208 3701 1290 3739
rect 1208 3667 1232 3701
rect 1266 3667 1290 3701
rect 1208 3629 1290 3667
rect 1208 3595 1232 3629
rect 1266 3595 1290 3629
rect 1208 3557 1290 3595
rect 1208 3523 1232 3557
rect 1266 3523 1290 3557
rect 1208 3485 1290 3523
rect 1208 3451 1232 3485
rect 1266 3451 1290 3485
rect 1208 3413 1290 3451
rect 1208 3379 1232 3413
rect 1266 3379 1290 3413
rect 1208 3341 1290 3379
rect 1208 3307 1232 3341
rect 1266 3307 1290 3341
rect 1208 3269 1290 3307
rect 1208 3235 1232 3269
rect 1266 3235 1290 3269
rect 1208 3197 1290 3235
rect 1208 3163 1232 3197
rect 1266 3163 1290 3197
rect 1208 3125 1290 3163
rect 1208 3091 1232 3125
rect 1266 3091 1290 3125
rect 1208 3053 1290 3091
rect 1208 3019 1232 3053
rect 1266 3019 1290 3053
rect 1208 2981 1290 3019
rect 1208 2947 1232 2981
rect 1266 2947 1290 2981
rect 1208 2909 1290 2947
rect 1208 2875 1232 2909
rect 1266 2875 1290 2909
rect 1208 2837 1290 2875
rect 1208 2803 1232 2837
rect 1266 2803 1290 2837
rect 1208 2765 1290 2803
rect 1208 2731 1232 2765
rect 1266 2731 1290 2765
rect 1208 2693 1290 2731
rect 1208 2659 1232 2693
rect 1266 2659 1290 2693
rect 1208 2621 1290 2659
rect 1208 2587 1232 2621
rect 1266 2587 1290 2621
rect 1208 2549 1290 2587
rect 1208 2515 1232 2549
rect 1266 2515 1290 2549
rect 1208 2477 1290 2515
rect 1208 2443 1232 2477
rect 1266 2443 1290 2477
rect 1208 2405 1290 2443
rect 1208 2371 1232 2405
rect 1266 2371 1290 2405
rect 1208 2333 1290 2371
rect 1208 2299 1232 2333
rect 1266 2299 1290 2333
rect 1208 2261 1290 2299
rect 1208 2227 1232 2261
rect 1266 2227 1290 2261
rect 1208 2189 1290 2227
rect 1208 2155 1232 2189
rect 1266 2155 1290 2189
rect 1208 2117 1290 2155
rect 1208 2083 1232 2117
rect 1266 2083 1290 2117
rect 1208 2045 1290 2083
rect 1208 2011 1232 2045
rect 1266 2011 1290 2045
rect 1208 1973 1290 2011
rect 1208 1939 1232 1973
rect 1266 1939 1290 1973
rect 1208 1901 1290 1939
rect 1208 1867 1232 1901
rect 1266 1867 1290 1901
rect 1208 1829 1290 1867
rect 1208 1795 1232 1829
rect 1266 1795 1290 1829
rect 1208 1757 1290 1795
rect 1208 1723 1232 1757
rect 1266 1723 1290 1757
rect 1208 1685 1290 1723
rect 1208 1651 1232 1685
rect 1266 1651 1290 1685
rect 1208 1613 1290 1651
rect 1208 1579 1232 1613
rect 1266 1579 1290 1613
rect 1208 1541 1290 1579
rect 1208 1507 1232 1541
rect 1266 1507 1290 1541
rect 1208 1469 1290 1507
rect 1208 1435 1232 1469
rect 1266 1435 1290 1469
rect 1208 1397 1290 1435
rect 1208 1363 1232 1397
rect 1266 1363 1290 1397
rect 1208 1325 1290 1363
rect 1208 1291 1232 1325
rect 1266 1291 1290 1325
rect 1208 1253 1290 1291
rect 1208 1219 1232 1253
rect 1266 1219 1290 1253
rect 1208 1181 1290 1219
rect 1208 1147 1232 1181
rect 1266 1147 1290 1181
rect 1208 1109 1290 1147
rect 1208 1075 1232 1109
rect 1266 1075 1290 1109
rect 1208 1037 1290 1075
rect 1208 1003 1232 1037
rect 1266 1003 1290 1037
rect 1208 965 1290 1003
rect 1208 931 1232 965
rect 1266 931 1290 965
rect 1208 893 1290 931
rect 1208 859 1232 893
rect 1266 859 1290 893
rect 1208 821 1290 859
rect 1208 787 1232 821
rect 1266 787 1290 821
rect 1208 749 1290 787
rect 1208 715 1232 749
rect 1266 715 1290 749
rect 1208 677 1290 715
rect 1208 643 1232 677
rect 1266 643 1290 677
rect 1208 605 1290 643
rect 1208 571 1232 605
rect 1266 571 1290 605
rect 1208 533 1290 571
rect 1208 499 1232 533
rect 1266 499 1290 533
rect 1208 461 1290 499
rect 1208 427 1232 461
rect 1266 427 1290 461
rect 1208 389 1290 427
rect 1208 355 1232 389
rect 1266 355 1290 389
rect 1208 317 1290 355
rect 1208 283 1232 317
rect 1266 283 1290 317
rect 1208 245 1290 283
rect 1208 211 1232 245
rect 1266 211 1290 245
rect 1208 173 1290 211
rect 1208 139 1232 173
rect 1266 139 1290 173
rect 1208 101 1290 139
rect 1208 67 1232 101
rect 1266 67 1290 101
rect 1208 29 1290 67
rect -1140 -43 -1058 -5
rect -1140 -77 -1116 -43
rect -1082 -77 -1058 -43
rect -1140 -115 -1058 -77
rect -1140 -149 -1116 -115
rect -1082 -149 -1058 -115
rect -1140 -187 -1058 -149
rect -1140 -221 -1116 -187
rect -1082 -221 -1058 -187
rect -1140 -259 -1058 -221
rect -1140 -293 -1116 -259
rect -1082 -293 -1058 -259
rect -1140 -331 -1058 -293
rect -1140 -365 -1116 -331
rect -1082 -365 -1058 -331
rect -1140 -403 -1058 -365
rect -1140 -437 -1116 -403
rect -1082 -437 -1058 -403
rect -1140 -475 -1058 -437
rect -1140 -509 -1116 -475
rect -1082 -509 -1058 -475
rect -1140 -547 -1058 -509
rect -1140 -581 -1116 -547
rect -1082 -581 -1058 -547
rect -1140 -619 -1058 -581
rect -1140 -653 -1116 -619
rect -1082 -653 -1058 -619
rect 1208 -5 1232 29
rect 1266 -5 1290 29
rect 1208 -43 1290 -5
rect 1208 -77 1232 -43
rect 1266 -77 1290 -43
rect 1208 -115 1290 -77
rect 1208 -149 1232 -115
rect 1266 -149 1290 -115
rect 1208 -187 1290 -149
rect 1208 -221 1232 -187
rect 1266 -221 1290 -187
rect 1208 -259 1290 -221
rect 1208 -293 1232 -259
rect 1266 -293 1290 -259
rect 1208 -331 1290 -293
rect 1208 -365 1232 -331
rect 1266 -365 1290 -331
rect 1208 -403 1290 -365
rect 1208 -437 1232 -403
rect 1266 -437 1290 -403
rect 1208 -475 1290 -437
rect 1208 -509 1232 -475
rect 1266 -509 1290 -475
rect 1208 -547 1290 -509
rect 1208 -581 1232 -547
rect 1266 -581 1290 -547
rect 1208 -619 1290 -581
rect -1140 -691 -1058 -653
rect -1140 -725 -1116 -691
rect -1082 -725 -1058 -691
rect -1140 -763 -1058 -725
rect -1140 -797 -1116 -763
rect -1082 -797 -1058 -763
rect -1140 -835 -1058 -797
rect -1140 -869 -1116 -835
rect -1082 -869 -1058 -835
rect -296 -650 460 -643
rect -296 -702 -289 -650
rect -237 -702 -215 -650
rect -163 -702 -141 -650
rect -89 -702 -67 -650
rect -15 -702 7 -650
rect 59 -702 81 -650
rect 133 -702 155 -650
rect 207 -702 229 -650
rect 281 -702 303 -650
rect 355 -702 377 -650
rect 429 -702 460 -650
rect -296 -724 460 -702
rect -296 -776 -289 -724
rect -237 -776 -215 -724
rect -163 -776 -141 -724
rect -89 -776 -67 -724
rect -15 -776 7 -724
rect 59 -776 81 -724
rect 133 -776 155 -724
rect 207 -776 229 -724
rect 281 -776 303 -724
rect 355 -776 377 -724
rect 429 -776 460 -724
rect -296 -798 460 -776
rect -296 -850 -289 -798
rect -237 -850 -215 -798
rect -163 -850 -141 -798
rect -89 -850 -67 -798
rect -15 -850 7 -798
rect 59 -850 81 -798
rect 133 -850 155 -798
rect 207 -850 229 -798
rect 281 -850 303 -798
rect 355 -850 377 -798
rect 429 -850 460 -798
rect -296 -857 460 -850
rect 1208 -653 1232 -619
rect 1266 -653 1290 -619
rect 1208 -691 1290 -653
rect 1208 -725 1232 -691
rect 1266 -725 1290 -691
rect 1208 -763 1290 -725
rect 1208 -797 1232 -763
rect 1266 -797 1290 -763
rect 1208 -835 1290 -797
rect -1140 -907 -1058 -869
rect -1140 -941 -1116 -907
rect -1082 -941 -1058 -907
rect -1140 -979 -1058 -941
rect -1140 -1013 -1116 -979
rect -1082 -1013 -1058 -979
rect -1140 -1051 -1058 -1013
rect -1140 -1085 -1116 -1051
rect -1082 -1085 -1058 -1051
rect -1140 -1100 -1058 -1085
rect 1208 -869 1232 -835
rect 1266 -869 1290 -835
rect 1208 -907 1290 -869
rect 1208 -941 1232 -907
rect 1266 -941 1290 -907
rect 1208 -979 1290 -941
rect 1208 -1013 1232 -979
rect 1266 -1013 1290 -979
rect 1208 -1051 1290 -1013
rect 1208 -1085 1232 -1051
rect 1266 -1085 1290 -1051
rect 1208 -1100 1290 -1085
rect -1140 -1124 1290 -1100
rect -1140 -1158 -988 -1124
rect -954 -1158 -916 -1124
rect -882 -1158 -844 -1124
rect -810 -1158 -772 -1124
rect -738 -1158 -700 -1124
rect -666 -1158 -628 -1124
rect -594 -1158 -556 -1124
rect -522 -1158 -484 -1124
rect -450 -1158 -412 -1124
rect -378 -1158 -340 -1124
rect -306 -1158 -268 -1124
rect -234 -1158 -196 -1124
rect -162 -1158 -124 -1124
rect -90 -1158 -52 -1124
rect -18 -1158 20 -1124
rect 54 -1158 92 -1124
rect 126 -1158 164 -1124
rect 198 -1158 236 -1124
rect 270 -1158 308 -1124
rect 342 -1158 380 -1124
rect 414 -1158 452 -1124
rect 486 -1158 524 -1124
rect 558 -1158 596 -1124
rect 630 -1158 668 -1124
rect 702 -1158 740 -1124
rect 774 -1158 812 -1124
rect 846 -1158 884 -1124
rect 918 -1158 956 -1124
rect 990 -1158 1028 -1124
rect 1062 -1158 1100 -1124
rect 1134 -1158 1290 -1124
rect -1140 -1182 1290 -1158
<< via1 >>
rect 17 5933 133 5939
rect 17 67 22 5933
rect 22 67 128 5933
rect 128 67 133 5933
rect 17 63 133 67
rect -289 -659 -237 -650
rect -289 -693 -280 -659
rect -280 -693 -246 -659
rect -246 -693 -237 -659
rect -289 -702 -237 -693
rect -215 -659 -163 -650
rect -215 -693 -206 -659
rect -206 -693 -172 -659
rect -172 -693 -163 -659
rect -215 -702 -163 -693
rect -141 -659 -89 -650
rect -141 -693 -132 -659
rect -132 -693 -98 -659
rect -98 -693 -89 -659
rect -141 -702 -89 -693
rect -67 -659 -15 -650
rect -67 -693 -58 -659
rect -58 -693 -24 -659
rect -24 -693 -15 -659
rect -67 -702 -15 -693
rect 7 -659 59 -650
rect 7 -693 16 -659
rect 16 -693 50 -659
rect 50 -693 59 -659
rect 7 -702 59 -693
rect 81 -659 133 -650
rect 81 -693 90 -659
rect 90 -693 124 -659
rect 124 -693 133 -659
rect 81 -702 133 -693
rect 155 -659 207 -650
rect 155 -693 164 -659
rect 164 -693 198 -659
rect 198 -693 207 -659
rect 155 -702 207 -693
rect 229 -659 281 -650
rect 229 -693 238 -659
rect 238 -693 272 -659
rect 272 -693 281 -659
rect 229 -702 281 -693
rect 303 -659 355 -650
rect 303 -693 312 -659
rect 312 -693 346 -659
rect 346 -693 355 -659
rect 303 -702 355 -693
rect 377 -659 429 -650
rect 377 -693 386 -659
rect 386 -693 420 -659
rect 420 -693 429 -659
rect 377 -702 429 -693
rect -289 -733 -237 -724
rect -289 -767 -280 -733
rect -280 -767 -246 -733
rect -246 -767 -237 -733
rect -289 -776 -237 -767
rect -215 -733 -163 -724
rect -215 -767 -206 -733
rect -206 -767 -172 -733
rect -172 -767 -163 -733
rect -215 -776 -163 -767
rect -141 -733 -89 -724
rect -141 -767 -132 -733
rect -132 -767 -98 -733
rect -98 -767 -89 -733
rect -141 -776 -89 -767
rect -67 -733 -15 -724
rect -67 -767 -58 -733
rect -58 -767 -24 -733
rect -24 -767 -15 -733
rect -67 -776 -15 -767
rect 7 -733 59 -724
rect 7 -767 16 -733
rect 16 -767 50 -733
rect 50 -767 59 -733
rect 7 -776 59 -767
rect 81 -733 133 -724
rect 81 -767 90 -733
rect 90 -767 124 -733
rect 124 -767 133 -733
rect 81 -776 133 -767
rect 155 -733 207 -724
rect 155 -767 164 -733
rect 164 -767 198 -733
rect 198 -767 207 -733
rect 155 -776 207 -767
rect 229 -733 281 -724
rect 229 -767 238 -733
rect 238 -767 272 -733
rect 272 -767 281 -733
rect 229 -776 281 -767
rect 303 -733 355 -724
rect 303 -767 312 -733
rect 312 -767 346 -733
rect 346 -767 355 -733
rect 303 -776 355 -767
rect 377 -733 429 -724
rect 377 -767 386 -733
rect 386 -767 420 -733
rect 420 -767 429 -733
rect 377 -776 429 -767
rect -289 -807 -237 -798
rect -289 -841 -280 -807
rect -280 -841 -246 -807
rect -246 -841 -237 -807
rect -289 -850 -237 -841
rect -215 -807 -163 -798
rect -215 -841 -206 -807
rect -206 -841 -172 -807
rect -172 -841 -163 -807
rect -215 -850 -163 -841
rect -141 -807 -89 -798
rect -141 -841 -132 -807
rect -132 -841 -98 -807
rect -98 -841 -89 -807
rect -141 -850 -89 -841
rect -67 -807 -15 -798
rect -67 -841 -58 -807
rect -58 -841 -24 -807
rect -24 -841 -15 -807
rect -67 -850 -15 -841
rect 7 -807 59 -798
rect 7 -841 16 -807
rect 16 -841 50 -807
rect 50 -841 59 -807
rect 7 -850 59 -841
rect 81 -807 133 -798
rect 81 -841 90 -807
rect 90 -841 124 -807
rect 124 -841 133 -807
rect 81 -850 133 -841
rect 155 -807 207 -798
rect 155 -841 164 -807
rect 164 -841 198 -807
rect 198 -841 207 -807
rect 155 -850 207 -841
rect 229 -807 281 -798
rect 229 -841 238 -807
rect 238 -841 272 -807
rect 272 -841 281 -807
rect 229 -850 281 -841
rect 303 -807 355 -798
rect 303 -841 312 -807
rect 312 -841 346 -807
rect 346 -841 355 -807
rect 303 -850 355 -841
rect 377 -807 429 -798
rect 377 -841 386 -807
rect 386 -841 420 -807
rect 420 -841 429 -807
rect 377 -850 429 -841
<< metal2 >>
rect 11 5939 139 5945
rect 11 63 17 5939
rect 133 63 139 5939
rect 11 57 139 63
rect -296 -650 460 -643
rect -296 -702 -289 -650
rect -237 -702 -215 -650
rect -163 -702 -141 -650
rect -89 -702 -67 -650
rect -15 -702 7 -650
rect 59 -702 81 -650
rect 133 -702 155 -650
rect 207 -702 229 -650
rect 281 -702 303 -650
rect 355 -702 377 -650
rect 429 -702 460 -650
rect -296 -724 460 -702
rect -296 -776 -289 -724
rect -237 -776 -215 -724
rect -163 -776 -141 -724
rect -89 -776 -67 -724
rect -15 -776 7 -724
rect 59 -776 81 -724
rect 133 -776 155 -724
rect 207 -776 229 -724
rect 281 -776 303 -724
rect 355 -776 377 -724
rect 429 -776 460 -724
rect -296 -798 460 -776
rect -296 -850 -289 -798
rect -237 -850 -215 -798
rect -163 -850 -141 -798
rect -89 -850 -67 -798
rect -15 -850 7 -798
rect 59 -850 81 -798
rect 133 -850 155 -798
rect 207 -850 229 -798
rect 281 -850 303 -798
rect 355 -850 377 -798
rect 429 -850 460 -798
rect -296 -857 460 -850
<< labels >>
flabel comment s -936 226 -936 226 0 FreeSans 1600 0 0 0 S
flabel comment s 1085 226 1085 226 0 FreeSans 1600 0 0 0 S
flabel comment s 79 206 79 206 0 FreeSans 1600 0 0 0 D
flabel locali s -296 -857 460 -853 0 FreeSans 400 0 0 0 G
port 2 nsew
flabel locali s 1156 7140 1290 7182 0 FreeSans 400 0 0 0 PSUB
port 3 nsew
flabel locali s 8 43 142 47 0 FreeSans 400 0 0 0 D
port 4 nsew
flabel locali s 1046 9 1112 13 0 FreeSans 400 0 0 0 S
port 5 nsew
flabel locali s -962 9 -896 13 0 FreeSans 400 0 0 0 S
port 5 nsew
<< properties >>
string GDS_END 7059886
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 6939182
<< end >>
