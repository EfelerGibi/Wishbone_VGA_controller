magic
tech sky130A
magscale 1 2
timestamp 1683767628
use sky130_fd_io__com_bus_hookup  sky130_fd_io__com_bus_hookup_0
timestamp 1683767628
transform 1 0 0 0 1 0
box 0 -142 15000 39451
use sky130_fd_io__pad_esd  sky130_fd_io__pad_esd_0
timestamp 1683767628
transform 1 0 0 0 1 0
box 960 18991 14040 34071
<< properties >>
string GDS_END 11194916
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 11194814
<< end >>
