magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< metal1 >>
rect 222 0 258 52140
rect 294 0 330 52140
rect 366 51429 402 51770
rect 366 50639 402 51271
rect 366 49849 402 50481
rect 366 49059 402 49691
rect 366 48269 402 48901
rect 366 47479 402 48111
rect 366 46689 402 47321
rect 366 45899 402 46531
rect 366 45109 402 45741
rect 366 44319 402 44951
rect 366 43529 402 44161
rect 366 42739 402 43371
rect 366 41949 402 42581
rect 366 41159 402 41791
rect 366 40369 402 41001
rect 366 39579 402 40211
rect 366 38789 402 39421
rect 366 37999 402 38631
rect 366 37209 402 37841
rect 366 36419 402 37051
rect 366 35629 402 36261
rect 366 34839 402 35471
rect 366 34049 402 34681
rect 366 33259 402 33891
rect 366 32469 402 33101
rect 366 31679 402 32311
rect 366 30889 402 31521
rect 366 30099 402 30731
rect 366 29309 402 29941
rect 366 28519 402 29151
rect 366 27729 402 28361
rect 366 26939 402 27571
rect 366 26149 402 26781
rect 366 25359 402 25991
rect 366 24569 402 25201
rect 366 23779 402 24411
rect 366 22989 402 23621
rect 366 22199 402 22831
rect 366 21409 402 22041
rect 366 20619 402 21251
rect 366 19829 402 20461
rect 366 19039 402 19671
rect 366 18249 402 18881
rect 366 17459 402 18091
rect 366 16669 402 17301
rect 366 15879 402 16511
rect 366 15089 402 15721
rect 366 14299 402 14931
rect 366 13509 402 14141
rect 366 12719 402 13351
rect 366 11929 402 12561
rect 366 11139 402 11771
rect 366 10349 402 10981
rect 366 9559 402 10191
rect 366 8769 402 9401
rect 366 7979 402 8611
rect 366 7189 402 7821
rect 366 6399 402 7031
rect 366 5609 402 6241
rect 366 4819 402 5451
rect 366 4029 402 4661
rect 366 3239 402 3871
rect 366 2449 402 3081
rect 366 1659 402 2291
rect 366 869 402 1501
rect 366 370 402 711
rect 438 0 474 52140
rect 510 0 546 52140
<< metal2 >>
rect 284 51939 340 51948
rect 284 51874 340 51883
rect 0 51673 624 51721
rect 330 51549 438 51625
rect 0 51453 624 51501
rect 330 51295 438 51405
rect 0 51199 624 51247
rect 330 51075 438 51151
rect 0 50979 624 51027
rect 0 50883 624 50931
rect 330 50759 438 50835
rect 0 50663 624 50711
rect 330 50505 438 50615
rect 0 50409 624 50457
rect 330 50285 438 50361
rect 0 50189 624 50237
rect 0 50093 624 50141
rect 330 49969 438 50045
rect 0 49873 624 49921
rect 330 49715 438 49825
rect 0 49619 624 49667
rect 330 49495 438 49571
rect 0 49399 624 49447
rect 0 49303 624 49351
rect 330 49179 438 49255
rect 0 49083 624 49131
rect 330 48925 438 49035
rect 0 48829 624 48877
rect 330 48705 438 48781
rect 0 48609 624 48657
rect 0 48513 624 48561
rect 330 48389 438 48465
rect 0 48293 624 48341
rect 330 48135 438 48245
rect 0 48039 624 48087
rect 330 47915 438 47991
rect 0 47819 624 47867
rect 0 47723 624 47771
rect 330 47599 438 47675
rect 0 47503 624 47551
rect 330 47345 438 47455
rect 0 47249 624 47297
rect 330 47125 438 47201
rect 0 47029 624 47077
rect 0 46933 624 46981
rect 330 46809 438 46885
rect 0 46713 624 46761
rect 330 46555 438 46665
rect 0 46459 624 46507
rect 330 46335 438 46411
rect 0 46239 624 46287
rect 0 46143 624 46191
rect 330 46019 438 46095
rect 0 45923 624 45971
rect 330 45765 438 45875
rect 0 45669 624 45717
rect 330 45545 438 45621
rect 0 45449 624 45497
rect 0 45353 624 45401
rect 330 45229 438 45305
rect 0 45133 624 45181
rect 330 44975 438 45085
rect 0 44879 624 44927
rect 330 44755 438 44831
rect 0 44659 624 44707
rect 0 44563 624 44611
rect 330 44439 438 44515
rect 0 44343 624 44391
rect 330 44185 438 44295
rect 0 44089 624 44137
rect 330 43965 438 44041
rect 0 43869 624 43917
rect 0 43773 624 43821
rect 330 43649 438 43725
rect 0 43553 624 43601
rect 330 43395 438 43505
rect 0 43299 624 43347
rect 330 43175 438 43251
rect 0 43079 624 43127
rect 0 42983 624 43031
rect 330 42859 438 42935
rect 0 42763 624 42811
rect 330 42605 438 42715
rect 0 42509 624 42557
rect 330 42385 438 42461
rect 0 42289 624 42337
rect 0 42193 624 42241
rect 330 42069 438 42145
rect 0 41973 624 42021
rect 330 41815 438 41925
rect 0 41719 624 41767
rect 330 41595 438 41671
rect 0 41499 624 41547
rect 0 41403 624 41451
rect 330 41279 438 41355
rect 0 41183 624 41231
rect 330 41025 438 41135
rect 0 40929 624 40977
rect 330 40805 438 40881
rect 0 40709 624 40757
rect 0 40613 624 40661
rect 330 40489 438 40565
rect 0 40393 624 40441
rect 330 40235 438 40345
rect 0 40139 624 40187
rect 330 40015 438 40091
rect 0 39919 624 39967
rect 0 39823 624 39871
rect 330 39699 438 39775
rect 0 39603 624 39651
rect 330 39445 438 39555
rect 0 39349 624 39397
rect 330 39225 438 39301
rect 0 39129 624 39177
rect 0 39033 624 39081
rect 330 38909 438 38985
rect 0 38813 624 38861
rect 330 38655 438 38765
rect 0 38559 624 38607
rect 330 38435 438 38511
rect 0 38339 624 38387
rect 0 38243 624 38291
rect 330 38119 438 38195
rect 0 38023 624 38071
rect 330 37865 438 37975
rect 0 37769 624 37817
rect 330 37645 438 37721
rect 0 37549 624 37597
rect 0 37453 624 37501
rect 330 37329 438 37405
rect 0 37233 624 37281
rect 330 37075 438 37185
rect 0 36979 624 37027
rect 330 36855 438 36931
rect 0 36759 624 36807
rect 0 36663 624 36711
rect 330 36539 438 36615
rect 0 36443 624 36491
rect 330 36285 438 36395
rect 0 36189 624 36237
rect 330 36065 438 36141
rect 0 35969 624 36017
rect 0 35873 624 35921
rect 330 35749 438 35825
rect 0 35653 624 35701
rect 330 35495 438 35605
rect 0 35399 624 35447
rect 330 35275 438 35351
rect 0 35179 624 35227
rect 0 35083 624 35131
rect 330 34959 438 35035
rect 0 34863 624 34911
rect 330 34705 438 34815
rect 0 34609 624 34657
rect 330 34485 438 34561
rect 0 34389 624 34437
rect 0 34293 624 34341
rect 330 34169 438 34245
rect 0 34073 624 34121
rect 330 33915 438 34025
rect 0 33819 624 33867
rect 330 33695 438 33771
rect 0 33599 624 33647
rect 0 33503 624 33551
rect 330 33379 438 33455
rect 0 33283 624 33331
rect 330 33125 438 33235
rect 0 33029 624 33077
rect 330 32905 438 32981
rect 0 32809 624 32857
rect 0 32713 624 32761
rect 330 32589 438 32665
rect 0 32493 624 32541
rect 330 32335 438 32445
rect 0 32239 624 32287
rect 330 32115 438 32191
rect 0 32019 624 32067
rect 0 31923 624 31971
rect 330 31799 438 31875
rect 0 31703 624 31751
rect 330 31545 438 31655
rect 0 31449 624 31497
rect 330 31325 438 31401
rect 0 31229 624 31277
rect 0 31133 624 31181
rect 330 31009 438 31085
rect 0 30913 624 30961
rect 330 30755 438 30865
rect 0 30659 624 30707
rect 330 30535 438 30611
rect 0 30439 624 30487
rect 0 30343 624 30391
rect 330 30219 438 30295
rect 0 30123 624 30171
rect 330 29965 438 30075
rect 0 29869 624 29917
rect 330 29745 438 29821
rect 0 29649 624 29697
rect 0 29553 624 29601
rect 330 29429 438 29505
rect 0 29333 624 29381
rect 330 29175 438 29285
rect 0 29079 624 29127
rect 330 28955 438 29031
rect 0 28859 624 28907
rect 0 28763 624 28811
rect 330 28639 438 28715
rect 0 28543 624 28591
rect 330 28385 438 28495
rect 0 28289 624 28337
rect 330 28165 438 28241
rect 0 28069 624 28117
rect 0 27973 624 28021
rect 330 27849 438 27925
rect 0 27753 624 27801
rect 330 27595 438 27705
rect 0 27499 624 27547
rect 330 27375 438 27451
rect 0 27279 624 27327
rect 0 27183 624 27231
rect 330 27059 438 27135
rect 0 26963 624 27011
rect 330 26805 438 26915
rect 0 26709 624 26757
rect 330 26585 438 26661
rect 0 26489 624 26537
rect 0 26393 624 26441
rect 330 26269 438 26345
rect 0 26173 624 26221
rect 330 26015 438 26125
rect 0 25919 624 25967
rect 330 25795 438 25871
rect 0 25699 624 25747
rect 0 25603 624 25651
rect 330 25479 438 25555
rect 0 25383 624 25431
rect 330 25225 438 25335
rect 0 25129 624 25177
rect 330 25005 438 25081
rect 0 24909 624 24957
rect 0 24813 624 24861
rect 330 24689 438 24765
rect 0 24593 624 24641
rect 330 24435 438 24545
rect 0 24339 624 24387
rect 330 24215 438 24291
rect 0 24119 624 24167
rect 0 24023 624 24071
rect 330 23899 438 23975
rect 0 23803 624 23851
rect 330 23645 438 23755
rect 0 23549 624 23597
rect 330 23425 438 23501
rect 0 23329 624 23377
rect 0 23233 624 23281
rect 330 23109 438 23185
rect 0 23013 624 23061
rect 330 22855 438 22965
rect 0 22759 624 22807
rect 330 22635 438 22711
rect 0 22539 624 22587
rect 0 22443 624 22491
rect 330 22319 438 22395
rect 0 22223 624 22271
rect 330 22065 438 22175
rect 0 21969 624 22017
rect 330 21845 438 21921
rect 0 21749 624 21797
rect 0 21653 624 21701
rect 330 21529 438 21605
rect 0 21433 624 21481
rect 330 21275 438 21385
rect 0 21179 624 21227
rect 330 21055 438 21131
rect 0 20959 624 21007
rect 0 20863 624 20911
rect 330 20739 438 20815
rect 0 20643 624 20691
rect 330 20485 438 20595
rect 0 20389 624 20437
rect 330 20265 438 20341
rect 0 20169 624 20217
rect 0 20073 624 20121
rect 330 19949 438 20025
rect 0 19853 624 19901
rect 330 19695 438 19805
rect 0 19599 624 19647
rect 330 19475 438 19551
rect 0 19379 624 19427
rect 0 19283 624 19331
rect 330 19159 438 19235
rect 0 19063 624 19111
rect 330 18905 438 19015
rect 0 18809 624 18857
rect 330 18685 438 18761
rect 0 18589 624 18637
rect 0 18493 624 18541
rect 330 18369 438 18445
rect 0 18273 624 18321
rect 330 18115 438 18225
rect 0 18019 624 18067
rect 330 17895 438 17971
rect 0 17799 624 17847
rect 0 17703 624 17751
rect 330 17579 438 17655
rect 0 17483 624 17531
rect 330 17325 438 17435
rect 0 17229 624 17277
rect 330 17105 438 17181
rect 0 17009 624 17057
rect 0 16913 624 16961
rect 330 16789 438 16865
rect 0 16693 624 16741
rect 330 16535 438 16645
rect 0 16439 624 16487
rect 330 16315 438 16391
rect 0 16219 624 16267
rect 0 16123 624 16171
rect 330 15999 438 16075
rect 0 15903 624 15951
rect 330 15745 438 15855
rect 0 15649 624 15697
rect 330 15525 438 15601
rect 0 15429 624 15477
rect 0 15333 624 15381
rect 330 15209 438 15285
rect 0 15113 624 15161
rect 330 14955 438 15065
rect 0 14859 624 14907
rect 330 14735 438 14811
rect 0 14639 624 14687
rect 0 14543 624 14591
rect 330 14419 438 14495
rect 0 14323 624 14371
rect 330 14165 438 14275
rect 0 14069 624 14117
rect 330 13945 438 14021
rect 0 13849 624 13897
rect 0 13753 624 13801
rect 330 13629 438 13705
rect 0 13533 624 13581
rect 330 13375 438 13485
rect 0 13279 624 13327
rect 330 13155 438 13231
rect 0 13059 624 13107
rect 0 12963 624 13011
rect 330 12839 438 12915
rect 0 12743 624 12791
rect 330 12585 438 12695
rect 0 12489 624 12537
rect 330 12365 438 12441
rect 0 12269 624 12317
rect 0 12173 624 12221
rect 330 12049 438 12125
rect 0 11953 624 12001
rect 330 11795 438 11905
rect 0 11699 624 11747
rect 330 11575 438 11651
rect 0 11479 624 11527
rect 0 11383 624 11431
rect 330 11259 438 11335
rect 0 11163 624 11211
rect 330 11005 438 11115
rect 0 10909 624 10957
rect 330 10785 438 10861
rect 0 10689 624 10737
rect 0 10593 624 10641
rect 330 10469 438 10545
rect 0 10373 624 10421
rect 330 10215 438 10325
rect 0 10119 624 10167
rect 330 9995 438 10071
rect 0 9899 624 9947
rect 0 9803 624 9851
rect 330 9679 438 9755
rect 0 9583 624 9631
rect 330 9425 438 9535
rect 0 9329 624 9377
rect 330 9205 438 9281
rect 0 9109 624 9157
rect 0 9013 624 9061
rect 330 8889 438 8965
rect 0 8793 624 8841
rect 330 8635 438 8745
rect 0 8539 624 8587
rect 330 8415 438 8491
rect 0 8319 624 8367
rect 0 8223 624 8271
rect 330 8099 438 8175
rect 0 8003 624 8051
rect 330 7845 438 7955
rect 0 7749 624 7797
rect 330 7625 438 7701
rect 0 7529 624 7577
rect 0 7433 624 7481
rect 330 7309 438 7385
rect 0 7213 624 7261
rect 330 7055 438 7165
rect 0 6959 624 7007
rect 330 6835 438 6911
rect 0 6739 624 6787
rect 0 6643 624 6691
rect 330 6519 438 6595
rect 0 6423 624 6471
rect 330 6265 438 6375
rect 0 6169 624 6217
rect 330 6045 438 6121
rect 0 5949 624 5997
rect 0 5853 624 5901
rect 330 5729 438 5805
rect 0 5633 624 5681
rect 330 5475 438 5585
rect 0 5379 624 5427
rect 330 5255 438 5331
rect 0 5159 624 5207
rect 0 5063 624 5111
rect 330 4939 438 5015
rect 0 4843 624 4891
rect 330 4685 438 4795
rect 0 4589 624 4637
rect 330 4465 438 4541
rect 0 4369 624 4417
rect 0 4273 624 4321
rect 330 4149 438 4225
rect 0 4053 624 4101
rect 330 3895 438 4005
rect 0 3799 624 3847
rect 330 3675 438 3751
rect 0 3579 624 3627
rect 0 3483 624 3531
rect 330 3359 438 3435
rect 0 3263 624 3311
rect 330 3105 438 3215
rect 0 3009 624 3057
rect 330 2885 438 2961
rect 0 2789 624 2837
rect 0 2693 624 2741
rect 330 2569 438 2645
rect 0 2473 624 2521
rect 330 2315 438 2425
rect 0 2219 624 2267
rect 330 2095 438 2171
rect 0 1999 624 2047
rect 0 1903 624 1951
rect 330 1779 438 1855
rect 0 1683 624 1731
rect 330 1525 438 1635
rect 0 1429 624 1477
rect 330 1305 438 1381
rect 0 1209 624 1257
rect 0 1113 624 1161
rect 330 989 438 1065
rect 0 893 624 941
rect 330 735 438 845
rect 0 639 624 687
rect 330 515 438 591
rect 0 419 624 467
rect 284 257 340 266
rect 284 192 340 201
<< via2 >>
rect 284 51883 340 51939
rect 284 201 340 257
<< metal3 >>
rect 263 51939 361 51960
rect 263 51883 284 51939
rect 340 51883 361 51939
rect 263 51862 361 51883
rect 263 257 361 278
rect 263 201 284 257
rect 340 201 361 257
rect 263 180 361 201
use contact_9  contact_9_0
timestamp 1683767628
transform 1 0 279 0 1 192
box 0 0 1 1
use contact_9  contact_9_1
timestamp 1683767628
transform 1 0 279 0 1 51874
box 0 0 1 1
use sky130_fd_bd_sram__openram_dp_cell_cap_col_1  sky130_fd_bd_sram__openram_dp_cell_cap_col_0
timestamp 1683767628
transform -1 0 624 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col_1  sky130_fd_bd_sram__openram_dp_cell_cap_col_1
timestamp 1683767628
transform -1 0 624 0 -1 52140
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_dummy_1  sky130_fd_bd_sram__openram_dp_cell_dummy_0
timestamp 1683767628
transform -1 0 624 0 1 51350
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_0
timestamp 1683767628
transform -1 0 624 0 1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_1
timestamp 1683767628
transform -1 0 624 0 -1 790
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_2
timestamp 1683767628
transform -1 0 624 0 1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_3
timestamp 1683767628
transform -1 0 624 0 -1 25280
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_4
timestamp 1683767628
transform -1 0 624 0 1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_5
timestamp 1683767628
transform -1 0 624 0 -1 24490
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_6
timestamp 1683767628
transform -1 0 624 0 1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_7
timestamp 1683767628
transform -1 0 624 0 -1 23700
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_8
timestamp 1683767628
transform -1 0 624 0 1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_9
timestamp 1683767628
transform -1 0 624 0 -1 22910
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_10
timestamp 1683767628
transform -1 0 624 0 1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_11
timestamp 1683767628
transform -1 0 624 0 -1 22120
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_12
timestamp 1683767628
transform -1 0 624 0 1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_13
timestamp 1683767628
transform -1 0 624 0 -1 21330
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_14
timestamp 1683767628
transform -1 0 624 0 1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_15
timestamp 1683767628
transform -1 0 624 0 -1 20540
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_16
timestamp 1683767628
transform -1 0 624 0 1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_17
timestamp 1683767628
transform -1 0 624 0 -1 19750
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_18
timestamp 1683767628
transform -1 0 624 0 1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_19
timestamp 1683767628
transform -1 0 624 0 -1 18960
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_20
timestamp 1683767628
transform -1 0 624 0 1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_21
timestamp 1683767628
transform -1 0 624 0 -1 18170
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_22
timestamp 1683767628
transform -1 0 624 0 1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_23
timestamp 1683767628
transform -1 0 624 0 -1 17380
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_24
timestamp 1683767628
transform -1 0 624 0 1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_25
timestamp 1683767628
transform -1 0 624 0 -1 16590
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_26
timestamp 1683767628
transform -1 0 624 0 1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_27
timestamp 1683767628
transform -1 0 624 0 -1 15800
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_28
timestamp 1683767628
transform -1 0 624 0 1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_29
timestamp 1683767628
transform -1 0 624 0 -1 15010
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_30
timestamp 1683767628
transform -1 0 624 0 1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_31
timestamp 1683767628
transform -1 0 624 0 -1 14220
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_32
timestamp 1683767628
transform -1 0 624 0 1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_33
timestamp 1683767628
transform -1 0 624 0 -1 13430
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_34
timestamp 1683767628
transform -1 0 624 0 1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_35
timestamp 1683767628
transform -1 0 624 0 -1 12640
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_36
timestamp 1683767628
transform -1 0 624 0 1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_37
timestamp 1683767628
transform -1 0 624 0 -1 11850
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_38
timestamp 1683767628
transform -1 0 624 0 1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_39
timestamp 1683767628
transform -1 0 624 0 -1 11060
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_40
timestamp 1683767628
transform -1 0 624 0 1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_41
timestamp 1683767628
transform -1 0 624 0 -1 10270
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_42
timestamp 1683767628
transform -1 0 624 0 1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_43
timestamp 1683767628
transform -1 0 624 0 -1 9480
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_44
timestamp 1683767628
transform -1 0 624 0 1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_45
timestamp 1683767628
transform -1 0 624 0 -1 8690
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_46
timestamp 1683767628
transform -1 0 624 0 1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_47
timestamp 1683767628
transform -1 0 624 0 -1 7900
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_48
timestamp 1683767628
transform -1 0 624 0 1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_49
timestamp 1683767628
transform -1 0 624 0 -1 7110
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_50
timestamp 1683767628
transform -1 0 624 0 1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_51
timestamp 1683767628
transform -1 0 624 0 -1 6320
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_52
timestamp 1683767628
transform -1 0 624 0 1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_53
timestamp 1683767628
transform -1 0 624 0 -1 5530
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_54
timestamp 1683767628
transform -1 0 624 0 1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_55
timestamp 1683767628
transform -1 0 624 0 -1 4740
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_56
timestamp 1683767628
transform -1 0 624 0 1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_57
timestamp 1683767628
transform -1 0 624 0 -1 3950
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_58
timestamp 1683767628
transform -1 0 624 0 1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_59
timestamp 1683767628
transform -1 0 624 0 -1 3160
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_60
timestamp 1683767628
transform -1 0 624 0 1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_61
timestamp 1683767628
transform -1 0 624 0 -1 2370
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_62
timestamp 1683767628
transform -1 0 624 0 1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_63
timestamp 1683767628
transform -1 0 624 0 -1 1580
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_64
timestamp 1683767628
transform -1 0 624 0 -1 51350
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_65
timestamp 1683767628
transform -1 0 624 0 1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_66
timestamp 1683767628
transform -1 0 624 0 -1 50560
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_67
timestamp 1683767628
transform -1 0 624 0 1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_68
timestamp 1683767628
transform -1 0 624 0 -1 49770
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_69
timestamp 1683767628
transform -1 0 624 0 1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_70
timestamp 1683767628
transform -1 0 624 0 -1 48980
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_71
timestamp 1683767628
transform -1 0 624 0 1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_72
timestamp 1683767628
transform -1 0 624 0 -1 48190
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_73
timestamp 1683767628
transform -1 0 624 0 1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_74
timestamp 1683767628
transform -1 0 624 0 -1 47400
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_75
timestamp 1683767628
transform -1 0 624 0 1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_76
timestamp 1683767628
transform -1 0 624 0 -1 46610
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_77
timestamp 1683767628
transform -1 0 624 0 1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_78
timestamp 1683767628
transform -1 0 624 0 -1 45820
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_79
timestamp 1683767628
transform -1 0 624 0 1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_80
timestamp 1683767628
transform -1 0 624 0 -1 45030
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_81
timestamp 1683767628
transform -1 0 624 0 1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_82
timestamp 1683767628
transform -1 0 624 0 -1 44240
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_83
timestamp 1683767628
transform -1 0 624 0 1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_84
timestamp 1683767628
transform -1 0 624 0 -1 43450
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_85
timestamp 1683767628
transform -1 0 624 0 1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_86
timestamp 1683767628
transform -1 0 624 0 -1 42660
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_87
timestamp 1683767628
transform -1 0 624 0 1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_88
timestamp 1683767628
transform -1 0 624 0 -1 41870
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_89
timestamp 1683767628
transform -1 0 624 0 1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_90
timestamp 1683767628
transform -1 0 624 0 -1 41080
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_91
timestamp 1683767628
transform -1 0 624 0 1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_92
timestamp 1683767628
transform -1 0 624 0 -1 40290
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_93
timestamp 1683767628
transform -1 0 624 0 1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_94
timestamp 1683767628
transform -1 0 624 0 -1 39500
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_95
timestamp 1683767628
transform -1 0 624 0 1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_96
timestamp 1683767628
transform -1 0 624 0 -1 38710
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_97
timestamp 1683767628
transform -1 0 624 0 1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_98
timestamp 1683767628
transform -1 0 624 0 -1 37920
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_99
timestamp 1683767628
transform -1 0 624 0 1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_100
timestamp 1683767628
transform -1 0 624 0 -1 37130
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_101
timestamp 1683767628
transform -1 0 624 0 1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_102
timestamp 1683767628
transform -1 0 624 0 -1 36340
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_103
timestamp 1683767628
transform -1 0 624 0 1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_104
timestamp 1683767628
transform -1 0 624 0 -1 35550
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_105
timestamp 1683767628
transform -1 0 624 0 1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_106
timestamp 1683767628
transform -1 0 624 0 -1 34760
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_107
timestamp 1683767628
transform -1 0 624 0 1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_108
timestamp 1683767628
transform -1 0 624 0 -1 33970
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_109
timestamp 1683767628
transform -1 0 624 0 1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_110
timestamp 1683767628
transform -1 0 624 0 -1 33180
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_111
timestamp 1683767628
transform -1 0 624 0 1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_112
timestamp 1683767628
transform -1 0 624 0 -1 32390
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_113
timestamp 1683767628
transform -1 0 624 0 1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_114
timestamp 1683767628
transform -1 0 624 0 -1 31600
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_115
timestamp 1683767628
transform -1 0 624 0 1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_116
timestamp 1683767628
transform -1 0 624 0 -1 30810
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_117
timestamp 1683767628
transform -1 0 624 0 1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_118
timestamp 1683767628
transform -1 0 624 0 -1 30020
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_119
timestamp 1683767628
transform -1 0 624 0 1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_120
timestamp 1683767628
transform -1 0 624 0 -1 29230
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_121
timestamp 1683767628
transform -1 0 624 0 1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_122
timestamp 1683767628
transform -1 0 624 0 -1 28440
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_123
timestamp 1683767628
transform -1 0 624 0 1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_124
timestamp 1683767628
transform -1 0 624 0 -1 27650
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_125
timestamp 1683767628
transform -1 0 624 0 1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_126
timestamp 1683767628
transform -1 0 624 0 -1 26860
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_127
timestamp 1683767628
transform -1 0 624 0 1 26070
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_replica_1  sky130_fd_bd_sram__openram_dp_cell_replica_128
timestamp 1683767628
transform -1 0 624 0 -1 26070
box -42 -105 650 421
<< labels >>
rlabel metal1 s 384 32930 384 32930 4 vdd
port 1 nsew
rlabel metal1 s 384 48730 384 48730 4 vdd
port 1 nsew
rlabel metal1 s 384 29479 384 29479 4 vdd
port 1 nsew
rlabel metal1 s 384 42909 384 42909 4 vdd
port 1 nsew
rlabel metal1 s 384 50019 384 50019 4 vdd
port 1 nsew
rlabel metal1 s 384 45279 384 45279 4 vdd
port 1 nsew
rlabel metal1 s 384 33720 384 33720 4 vdd
port 1 nsew
rlabel metal1 s 384 36589 384 36589 4 vdd
port 1 nsew
rlabel metal1 s 384 26610 384 26610 4 vdd
port 1 nsew
rlabel metal1 s 384 51599 384 51599 4 vdd
port 1 nsew
rlabel metal1 s 384 28190 384 28190 4 vdd
port 1 nsew
rlabel metal1 s 384 51100 384 51100 4 vdd
port 1 nsew
rlabel metal1 s 384 38169 384 38169 4 vdd
port 1 nsew
rlabel metal1 s 384 32639 384 32639 4 vdd
port 1 nsew
rlabel metal1 s 384 49520 384 49520 4 vdd
port 1 nsew
rlabel metal1 s 384 38959 384 38959 4 vdd
port 1 nsew
rlabel metal1 s 384 41620 384 41620 4 vdd
port 1 nsew
rlabel metal1 s 384 43990 384 43990 4 vdd
port 1 nsew
rlabel metal1 s 384 34510 384 34510 4 vdd
port 1 nsew
rlabel metal1 s 384 37670 384 37670 4 vdd
port 1 nsew
rlabel metal1 s 384 31849 384 31849 4 vdd
port 1 nsew
rlabel metal1 s 384 43699 384 43699 4 vdd
port 1 nsew
rlabel metal1 s 384 29770 384 29770 4 vdd
port 1 nsew
rlabel metal1 s 384 33429 384 33429 4 vdd
port 1 nsew
rlabel metal1 s 384 28689 384 28689 4 vdd
port 1 nsew
rlabel metal1 s 384 40539 384 40539 4 vdd
port 1 nsew
rlabel metal1 s 384 40040 384 40040 4 vdd
port 1 nsew
rlabel metal1 s 384 27400 384 27400 4 vdd
port 1 nsew
rlabel metal1 s 384 46360 384 46360 4 vdd
port 1 nsew
rlabel metal1 s 384 34219 384 34219 4 vdd
port 1 nsew
rlabel metal1 s 384 46069 384 46069 4 vdd
port 1 nsew
rlabel metal1 s 384 26319 384 26319 4 vdd
port 1 nsew
rlabel metal1 s 384 50809 384 50809 4 vdd
port 1 nsew
rlabel metal1 s 384 47150 384 47150 4 vdd
port 1 nsew
rlabel metal1 s 384 49229 384 49229 4 vdd
port 1 nsew
rlabel metal1 s 384 46859 384 46859 4 vdd
port 1 nsew
rlabel metal1 s 384 27109 384 27109 4 vdd
port 1 nsew
rlabel metal1 s 384 47649 384 47649 4 vdd
port 1 nsew
rlabel metal1 s 384 44780 384 44780 4 vdd
port 1 nsew
rlabel metal1 s 384 31059 384 31059 4 vdd
port 1 nsew
rlabel metal1 s 384 28980 384 28980 4 vdd
port 1 nsew
rlabel metal1 s 384 44489 384 44489 4 vdd
port 1 nsew
rlabel metal1 s 384 38460 384 38460 4 vdd
port 1 nsew
rlabel metal1 s 384 30269 384 30269 4 vdd
port 1 nsew
rlabel metal1 s 384 36880 384 36880 4 vdd
port 1 nsew
rlabel metal1 s 384 31350 384 31350 4 vdd
port 1 nsew
rlabel metal1 s 384 40830 384 40830 4 vdd
port 1 nsew
rlabel metal1 s 384 42410 384 42410 4 vdd
port 1 nsew
rlabel metal1 s 384 48439 384 48439 4 vdd
port 1 nsew
rlabel metal1 s 384 32140 384 32140 4 vdd
port 1 nsew
rlabel metal1 s 384 43200 384 43200 4 vdd
port 1 nsew
rlabel metal1 s 384 47940 384 47940 4 vdd
port 1 nsew
rlabel metal1 s 384 42119 384 42119 4 vdd
port 1 nsew
rlabel metal1 s 384 35009 384 35009 4 vdd
port 1 nsew
rlabel metal1 s 384 35799 384 35799 4 vdd
port 1 nsew
rlabel metal1 s 384 39749 384 39749 4 vdd
port 1 nsew
rlabel metal1 s 384 30560 384 30560 4 vdd
port 1 nsew
rlabel metal1 s 384 36090 384 36090 4 vdd
port 1 nsew
rlabel metal1 s 384 50310 384 50310 4 vdd
port 1 nsew
rlabel metal1 s 384 37379 384 37379 4 vdd
port 1 nsew
rlabel metal1 s 384 41329 384 41329 4 vdd
port 1 nsew
rlabel metal1 s 384 35300 384 35300 4 vdd
port 1 nsew
rlabel metal1 s 384 45570 384 45570 4 vdd
port 1 nsew
rlabel metal1 s 384 27899 384 27899 4 vdd
port 1 nsew
rlabel metal1 s 384 39250 384 39250 4 vdd
port 1 nsew
rlabel metal1 s 240 26070 240 26070 4 br1
port 1067 nsew
rlabel metal1 s 384 15259 384 15259 4 vdd
port 1 nsew
rlabel metal1 s 384 19500 384 19500 4 vdd
port 1 nsew
rlabel metal1 s 384 8939 384 8939 4 vdd
port 1 nsew
rlabel metal1 s 384 10519 384 10519 4 vdd
port 1 nsew
rlabel metal1 s 384 12889 384 12889 4 vdd
port 1 nsew
rlabel metal1 s 384 17920 384 17920 4 vdd
port 1 nsew
rlabel metal1 s 384 25529 384 25529 4 vdd
port 1 nsew
rlabel metal1 s 384 2619 384 2619 4 vdd
port 1 nsew
rlabel metal1 s 384 23159 384 23159 4 vdd
port 1 nsew
rlabel metal1 s 384 13180 384 13180 4 vdd
port 1 nsew
rlabel metal1 s 384 6569 384 6569 4 vdd
port 1 nsew
rlabel metal1 s 384 3409 384 3409 4 vdd
port 1 nsew
rlabel metal1 s 384 24240 384 24240 4 vdd
port 1 nsew
rlabel metal1 s 384 9729 384 9729 4 vdd
port 1 nsew
rlabel metal1 s 384 4199 384 4199 4 vdd
port 1 nsew
rlabel metal1 s 384 23450 384 23450 4 vdd
port 1 nsew
rlabel metal1 s 384 14469 384 14469 4 vdd
port 1 nsew
rlabel metal1 s 384 22660 384 22660 4 vdd
port 1 nsew
rlabel metal1 s 384 9230 384 9230 4 vdd
port 1 nsew
rlabel metal1 s 384 10020 384 10020 4 vdd
port 1 nsew
rlabel metal1 s 384 11600 384 11600 4 vdd
port 1 nsew
rlabel metal1 s 384 21080 384 21080 4 vdd
port 1 nsew
rlabel metal1 s 384 4490 384 4490 4 vdd
port 1 nsew
rlabel metal1 s 384 18710 384 18710 4 vdd
port 1 nsew
rlabel metal1 s 384 21579 384 21579 4 vdd
port 1 nsew
rlabel metal1 s 384 3700 384 3700 4 vdd
port 1 nsew
rlabel metal1 s 384 23949 384 23949 4 vdd
port 1 nsew
rlabel metal1 s 384 25820 384 25820 4 vdd
port 1 nsew
rlabel metal1 s 384 24739 384 24739 4 vdd
port 1 nsew
rlabel metal1 s 384 14760 384 14760 4 vdd
port 1 nsew
rlabel metal1 s 384 21870 384 21870 4 vdd
port 1 nsew
rlabel metal1 s 384 13970 384 13970 4 vdd
port 1 nsew
rlabel metal1 s 384 10810 384 10810 4 vdd
port 1 nsew
rlabel metal1 s 384 19999 384 19999 4 vdd
port 1 nsew
rlabel metal1 s 384 2910 384 2910 4 vdd
port 1 nsew
rlabel metal1 s 384 20290 384 20290 4 vdd
port 1 nsew
rlabel metal1 s 384 1829 384 1829 4 vdd
port 1 nsew
rlabel metal1 s 384 22369 384 22369 4 vdd
port 1 nsew
rlabel metal1 s 384 11309 384 11309 4 vdd
port 1 nsew
rlabel metal1 s 384 16839 384 16839 4 vdd
port 1 nsew
rlabel metal1 s 384 17629 384 17629 4 vdd
port 1 nsew
rlabel metal1 s 384 4989 384 4989 4 vdd
port 1 nsew
rlabel metal1 s 384 20789 384 20789 4 vdd
port 1 nsew
rlabel metal1 s 384 7359 384 7359 4 vdd
port 1 nsew
rlabel metal1 s 384 19209 384 19209 4 vdd
port 1 nsew
rlabel metal1 s 384 8149 384 8149 4 vdd
port 1 nsew
rlabel metal1 s 384 15550 384 15550 4 vdd
port 1 nsew
rlabel metal1 s 384 1039 384 1039 4 vdd
port 1 nsew
rlabel metal1 s 384 17130 384 17130 4 vdd
port 1 nsew
rlabel metal1 s 384 13679 384 13679 4 vdd
port 1 nsew
rlabel metal1 s 384 5779 384 5779 4 vdd
port 1 nsew
rlabel metal1 s 384 18419 384 18419 4 vdd
port 1 nsew
rlabel metal1 s 384 1330 384 1330 4 vdd
port 1 nsew
rlabel metal1 s 384 6070 384 6070 4 vdd
port 1 nsew
rlabel metal1 s 384 16049 384 16049 4 vdd
port 1 nsew
rlabel metal1 s 384 16340 384 16340 4 vdd
port 1 nsew
rlabel metal1 s 384 2120 384 2120 4 vdd
port 1 nsew
rlabel metal1 s 384 5280 384 5280 4 vdd
port 1 nsew
rlabel metal1 s 384 12390 384 12390 4 vdd
port 1 nsew
rlabel metal1 s 384 7650 384 7650 4 vdd
port 1 nsew
rlabel metal1 s 384 6860 384 6860 4 vdd
port 1 nsew
rlabel metal1 s 384 540 384 540 4 vdd
port 1 nsew
rlabel metal1 s 384 12099 384 12099 4 vdd
port 1 nsew
rlabel metal1 s 384 25030 384 25030 4 vdd
port 1 nsew
rlabel metal1 s 312 26070 312 26070 4 bl1
port 1068 nsew
rlabel metal1 s 384 8440 384 8440 4 vdd
port 1 nsew
rlabel metal1 s 528 26070 528 26070 4 bl0
port 804 nsew
rlabel metal1 s 456 26070 456 26070 4 br0
port 806 nsew
rlabel metal2 s 384 26623 384 26623 4 gnd
port 2 nsew
rlabel metal2 s 384 47400 384 47400 4 gnd
port 2 nsew
rlabel metal2 s 384 35313 384 35313 4 gnd
port 2 nsew
rlabel metal2 s 384 35787 384 35787 4 gnd
port 2 nsew
rlabel metal2 s 384 29230 384 29230 4 gnd
port 2 nsew
rlabel metal2 s 384 42107 384 42107 4 gnd
port 2 nsew
rlabel metal2 s 384 31047 384 31047 4 gnd
port 2 nsew
rlabel metal2 s 384 38947 384 38947 4 gnd
port 2 nsew
rlabel metal2 s 384 28677 384 28677 4 gnd
port 2 nsew
rlabel metal2 s 384 41870 384 41870 4 gnd
port 2 nsew
rlabel metal2 s 384 49770 384 49770 4 gnd
port 2 nsew
rlabel metal2 s 384 31363 384 31363 4 gnd
port 2 nsew
rlabel metal2 s 384 45820 384 45820 4 gnd
port 2 nsew
rlabel metal2 s 384 32153 384 32153 4 gnd
port 2 nsew
rlabel metal2 s 384 50797 384 50797 4 gnd
port 2 nsew
rlabel metal2 s 384 36577 384 36577 4 gnd
port 2 nsew
rlabel metal2 s 384 38157 384 38157 4 gnd
port 2 nsew
rlabel metal2 s 384 47163 384 47163 4 gnd
port 2 nsew
rlabel metal2 s 384 36893 384 36893 4 gnd
port 2 nsew
rlabel metal2 s 384 32627 384 32627 4 gnd
port 2 nsew
rlabel metal2 s 384 38710 384 38710 4 gnd
port 2 nsew
rlabel metal2 s 384 32390 384 32390 4 gnd
port 2 nsew
rlabel metal2 s 384 34760 384 34760 4 gnd
port 2 nsew
rlabel metal2 s 384 44003 384 44003 4 gnd
port 2 nsew
rlabel metal2 s 384 50560 384 50560 4 gnd
port 2 nsew
rlabel metal2 s 384 36103 384 36103 4 gnd
port 2 nsew
rlabel metal2 s 384 42897 384 42897 4 gnd
port 2 nsew
rlabel metal2 s 384 40527 384 40527 4 gnd
port 2 nsew
rlabel metal2 s 384 37130 384 37130 4 gnd
port 2 nsew
rlabel metal2 s 384 45030 384 45030 4 gnd
port 2 nsew
rlabel metal2 s 384 28993 384 28993 4 gnd
port 2 nsew
rlabel metal2 s 384 43213 384 43213 4 gnd
port 2 nsew
rlabel metal2 s 384 33417 384 33417 4 gnd
port 2 nsew
rlabel metal2 s 384 46373 384 46373 4 gnd
port 2 nsew
rlabel metal2 s 384 26860 384 26860 4 gnd
port 2 nsew
rlabel metal2 s 384 40843 384 40843 4 gnd
port 2 nsew
rlabel metal2 s 384 30257 384 30257 4 gnd
port 2 nsew
rlabel metal2 s 384 43687 384 43687 4 gnd
port 2 nsew
rlabel metal2 s 384 41317 384 41317 4 gnd
port 2 nsew
rlabel metal2 s 384 41080 384 41080 4 gnd
port 2 nsew
rlabel metal2 s 384 27887 384 27887 4 gnd
port 2 nsew
rlabel metal2 s 384 38473 384 38473 4 gnd
port 2 nsew
rlabel metal2 s 384 30020 384 30020 4 gnd
port 2 nsew
rlabel metal2 s 384 33970 384 33970 4 gnd
port 2 nsew
rlabel metal2 s 384 33180 384 33180 4 gnd
port 2 nsew
rlabel metal2 s 384 40290 384 40290 4 gnd
port 2 nsew
rlabel metal2 s 384 44793 384 44793 4 gnd
port 2 nsew
rlabel metal2 s 384 31600 384 31600 4 gnd
port 2 nsew
rlabel metal2 s 384 28440 384 28440 4 gnd
port 2 nsew
rlabel metal2 s 384 36340 384 36340 4 gnd
port 2 nsew
rlabel metal2 s 384 30810 384 30810 4 gnd
port 2 nsew
rlabel metal2 s 384 47953 384 47953 4 gnd
port 2 nsew
rlabel metal2 s 384 42423 384 42423 4 gnd
port 2 nsew
rlabel metal2 s 384 37683 384 37683 4 gnd
port 2 nsew
rlabel metal2 s 384 48190 384 48190 4 gnd
port 2 nsew
rlabel metal2 s 384 29467 384 29467 4 gnd
port 2 nsew
rlabel metal2 s 384 33733 384 33733 4 gnd
port 2 nsew
rlabel metal2 s 384 50007 384 50007 4 gnd
port 2 nsew
rlabel metal2 s 384 29783 384 29783 4 gnd
port 2 nsew
rlabel metal2 s 384 46057 384 46057 4 gnd
port 2 nsew
rlabel metal2 s 384 46847 384 46847 4 gnd
port 2 nsew
rlabel metal2 s 384 46610 384 46610 4 gnd
port 2 nsew
rlabel metal2 s 384 27097 384 27097 4 gnd
port 2 nsew
rlabel metal2 s 384 30573 384 30573 4 gnd
port 2 nsew
rlabel metal2 s 384 32943 384 32943 4 gnd
port 2 nsew
rlabel metal2 s 384 44477 384 44477 4 gnd
port 2 nsew
rlabel metal2 s 384 40053 384 40053 4 gnd
port 2 nsew
rlabel metal2 s 384 27650 384 27650 4 gnd
port 2 nsew
rlabel metal2 s 384 51113 384 51113 4 gnd
port 2 nsew
rlabel metal2 s 384 45583 384 45583 4 gnd
port 2 nsew
rlabel metal2 s 384 39500 384 39500 4 gnd
port 2 nsew
rlabel metal2 s 384 27413 384 27413 4 gnd
port 2 nsew
rlabel metal2 s 384 45267 384 45267 4 gnd
port 2 nsew
rlabel metal2 s 384 28203 384 28203 4 gnd
port 2 nsew
rlabel metal2 s 384 39263 384 39263 4 gnd
port 2 nsew
rlabel metal2 s 384 48427 384 48427 4 gnd
port 2 nsew
rlabel metal2 s 384 49533 384 49533 4 gnd
port 2 nsew
rlabel metal2 s 384 41633 384 41633 4 gnd
port 2 nsew
rlabel metal2 s 384 26307 384 26307 4 gnd
port 2 nsew
rlabel metal2 s 384 39737 384 39737 4 gnd
port 2 nsew
rlabel metal2 s 384 34997 384 34997 4 gnd
port 2 nsew
rlabel metal2 s 384 51587 384 51587 4 gnd
port 2 nsew
rlabel metal2 s 384 37367 384 37367 4 gnd
port 2 nsew
rlabel metal2 s 384 49217 384 49217 4 gnd
port 2 nsew
rlabel metal2 s 384 47637 384 47637 4 gnd
port 2 nsew
rlabel metal2 s 384 48743 384 48743 4 gnd
port 2 nsew
rlabel metal2 s 384 31837 384 31837 4 gnd
port 2 nsew
rlabel metal2 s 384 34207 384 34207 4 gnd
port 2 nsew
rlabel metal2 s 384 48980 384 48980 4 gnd
port 2 nsew
rlabel metal2 s 384 51350 384 51350 4 gnd
port 2 nsew
rlabel metal2 s 384 42660 384 42660 4 gnd
port 2 nsew
rlabel metal2 s 384 37920 384 37920 4 gnd
port 2 nsew
rlabel metal2 s 384 34523 384 34523 4 gnd
port 2 nsew
rlabel metal2 s 384 35550 384 35550 4 gnd
port 2 nsew
rlabel metal2 s 384 50323 384 50323 4 gnd
port 2 nsew
rlabel metal2 s 384 44240 384 44240 4 gnd
port 2 nsew
rlabel metal2 s 384 43450 384 43450 4 gnd
port 2 nsew
rlabel metal2 s 312 51477 312 51477 4 wl1_130
port 1066 nsew
rlabel metal2 s 312 48063 312 48063 4 wl1_121
port 1048 nsew
rlabel metal2 s 312 43577 312 43577 4 wl1_110
port 1026 nsew
rlabel metal2 s 312 49643 312 49643 4 wl1_125
port 1056 nsew
rlabel metal2 s 312 44113 312 44113 4 wl1_111
port 1028 nsew
rlabel metal2 s 312 41743 312 41743 4 wl1_105
port 1016 nsew
rlabel metal2 s 312 44903 312 44903 4 wl1_113
port 1032 nsew
rlabel metal2 s 312 49107 312 49107 4 wl1_124
port 1054 nsew
rlabel metal2 s 312 42313 312 42313 4 wl0_107
port 1019 nsew
rlabel metal2 s 312 50433 312 50433 4 wl1_127
port 1060 nsew
rlabel metal2 s 312 49327 312 49327 4 wl0_124
port 1053 nsew
rlabel metal2 s 312 43007 312 43007 4 wl0_108
port 1021 nsew
rlabel metal2 s 312 50117 312 50117 4 wl0_126
port 1057 nsew
rlabel metal2 s 312 40637 312 40637 4 wl0_102
port 1009 nsew
rlabel metal2 s 312 45377 312 45377 4 wl0_114
port 1033 nsew
rlabel metal2 s 312 42533 312 42533 4 wl1_107
port 1020 nsew
rlabel metal2 s 312 48853 312 48853 4 wl1_123
port 1052 nsew
rlabel metal2 s 312 40417 312 40417 4 wl1_102
port 1010 nsew
rlabel metal2 s 312 47843 312 47843 4 wl0_121
port 1047 nsew
rlabel metal2 s 312 40953 312 40953 4 wl1_103
port 1012 nsew
rlabel metal2 s 312 46263 312 46263 4 wl0_117
port 1039 nsew
rlabel metal2 s 312 48537 312 48537 4 wl0_122
port 1049 nsew
rlabel metal2 s 312 39057 312 39057 4 wl0_98
port 1001 nsew
rlabel metal2 s 312 47747 312 47747 4 wl0_120
port 1045 nsew
rlabel metal2 s 312 39847 312 39847 4 wl0_100
port 1005 nsew
rlabel metal2 s 312 44683 312 44683 4 wl0_113
port 1031 nsew
rlabel metal2 s 312 42787 312 42787 4 wl1_108
port 1022 nsew
rlabel metal2 s 312 50687 312 50687 4 wl1_128
port 1062 nsew
rlabel metal2 s 312 47273 312 47273 4 wl1_119
port 1044 nsew
rlabel metal2 s 312 39627 312 39627 4 wl1_100
port 1006 nsew
rlabel metal2 s 312 43893 312 43893 4 wl0_111
port 1027 nsew
rlabel metal2 s 312 45947 312 45947 4 wl1_116
port 1038 nsew
rlabel metal2 s 312 39153 312 39153 4 wl0_99
port 1003 nsew
rlabel metal2 s 312 51223 312 51223 4 wl1_129
port 1064 nsew
rlabel metal2 s 312 46957 312 46957 4 wl0_118
port 1041 nsew
rlabel metal2 s 312 41523 312 41523 4 wl0_105
port 1015 nsew
rlabel metal2 s 312 43797 312 43797 4 wl0_110
port 1025 nsew
rlabel metal2 s 312 45157 312 45157 4 wl1_114
port 1034 nsew
rlabel metal2 s 312 44367 312 44367 4 wl1_112
port 1030 nsew
rlabel metal2 s 312 51697 312 51697 4 wl0_130
port 1065 nsew
rlabel metal2 s 312 45473 312 45473 4 wl0_115
port 1035 nsew
rlabel metal2 s 312 41997 312 41997 4 wl1_106
port 1018 nsew
rlabel metal2 s 312 48317 312 48317 4 wl1_122
port 1050 nsew
rlabel metal2 s 312 51003 312 51003 4 wl0_129
port 1063 nsew
rlabel metal2 s 312 40163 312 40163 4 wl1_101
port 1008 nsew
rlabel metal2 s 312 50213 312 50213 4 wl0_127
port 1059 nsew
rlabel metal2 s 312 50907 312 50907 4 wl0_128
port 1061 nsew
rlabel metal2 s 312 43103 312 43103 4 wl0_109
port 1023 nsew
rlabel metal2 s 312 45693 312 45693 4 wl1_115
port 1036 nsew
rlabel metal2 s 312 46167 312 46167 4 wl0_116
port 1037 nsew
rlabel metal2 s 312 46483 312 46483 4 wl1_117
port 1040 nsew
rlabel metal2 s 312 46737 312 46737 4 wl1_118
port 1042 nsew
rlabel metal2 s 312 39943 312 39943 4 wl0_101
port 1007 nsew
rlabel metal2 s 312 47527 312 47527 4 wl1_120
port 1046 nsew
rlabel metal2 s 312 40733 312 40733 4 wl0_103
port 1011 nsew
rlabel metal2 s 312 41427 312 41427 4 wl0_104
port 1013 nsew
rlabel metal2 s 312 39373 312 39373 4 wl1_99
port 1004 nsew
rlabel metal2 s 312 47053 312 47053 4 wl0_119
port 1043 nsew
rlabel metal2 s 312 49897 312 49897 4 wl1_126
port 1058 nsew
rlabel metal2 s 312 44587 312 44587 4 wl0_112
port 1029 nsew
rlabel metal2 s 312 42217 312 42217 4 wl0_106
port 1017 nsew
rlabel metal2 s 312 49423 312 49423 4 wl0_125
port 1055 nsew
rlabel metal2 s 312 48633 312 48633 4 wl0_123
port 1051 nsew
rlabel metal2 s 312 43323 312 43323 4 wl1_109
port 1024 nsew
rlabel metal2 s 312 41207 312 41207 4 wl1_104
port 1014 nsew
rlabel metal2 s 312 35107 312 35107 4 wl0_88
port 981 nsew
rlabel metal2 s 312 27207 312 27207 4 wl0_68
port 941 nsew
rlabel metal2 s 312 30683 312 30683 4 wl1_77
port 960 nsew
rlabel metal2 s 312 28787 312 28787 4 wl0_72
port 949 nsew
rlabel metal2 s 312 35677 312 35677 4 wl1_90
port 986 nsew
rlabel metal2 s 312 31157 312 31157 4 wl0_78
port 961 nsew
rlabel metal2 s 312 36687 312 36687 4 wl0_92
port 989 nsew
rlabel metal2 s 312 26513 312 26513 4 wl0_67
port 939 nsew
rlabel metal2 s 312 38837 312 38837 4 wl1_98
port 1002 nsew
rlabel metal2 s 312 36783 312 36783 4 wl0_93
port 991 nsew
rlabel metal2 s 312 33307 312 33307 4 wl1_84
port 974 nsew
rlabel metal2 s 312 30463 312 30463 4 wl0_77
port 959 nsew
rlabel metal2 s 312 29673 312 29673 4 wl0_75
port 955 nsew
rlabel metal2 s 312 31947 312 31947 4 wl0_80
port 965 nsew
rlabel metal2 s 312 36467 312 36467 4 wl1_92
port 990 nsew
rlabel metal2 s 312 32043 312 32043 4 wl0_81
port 967 nsew
rlabel metal2 s 312 31253 312 31253 4 wl0_79
port 963 nsew
rlabel metal2 s 312 38583 312 38583 4 wl1_97
port 1000 nsew
rlabel metal2 s 312 26197 312 26197 4 wl1_66
port 938 nsew
rlabel metal2 s 312 37257 312 37257 4 wl1_94
port 994 nsew
rlabel metal2 s 312 36213 312 36213 4 wl1_91
port 988 nsew
rlabel metal2 s 312 29103 312 29103 4 wl1_73
port 952 nsew
rlabel metal2 s 312 34413 312 34413 4 wl0_87
port 979 nsew
rlabel metal2 s 312 31473 312 31473 4 wl1_79
port 964 nsew
rlabel metal2 s 312 27997 312 27997 4 wl0_70
port 945 nsew
rlabel metal2 s 312 32263 312 32263 4 wl1_81
port 968 nsew
rlabel metal2 s 312 26733 312 26733 4 wl1_67
port 940 nsew
rlabel metal2 s 312 27777 312 27777 4 wl1_70
port 946 nsew
rlabel metal2 s 312 37477 312 37477 4 wl0_94
port 993 nsew
rlabel metal2 s 312 30367 312 30367 4 wl0_76
port 957 nsew
rlabel metal2 s 312 28883 312 28883 4 wl0_73
port 951 nsew
rlabel metal2 s 312 32833 312 32833 4 wl0_83
port 971 nsew
rlabel metal2 s 312 28313 312 28313 4 wl1_71
port 948 nsew
rlabel metal2 s 312 38363 312 38363 4 wl0_97
port 999 nsew
rlabel metal2 s 312 35897 312 35897 4 wl0_90
port 985 nsew
rlabel metal2 s 312 33843 312 33843 4 wl1_85
port 976 nsew
rlabel metal2 s 312 26987 312 26987 4 wl1_68
port 942 nsew
rlabel metal2 s 312 33053 312 33053 4 wl1_83
port 972 nsew
rlabel metal2 s 312 32517 312 32517 4 wl1_82
port 970 nsew
rlabel metal2 s 312 31727 312 31727 4 wl1_80
port 966 nsew
rlabel metal2 s 312 35423 312 35423 4 wl1_89
port 984 nsew
rlabel metal2 s 312 38267 312 38267 4 wl0_96
port 997 nsew
rlabel metal2 s 312 35993 312 35993 4 wl0_91
port 987 nsew
rlabel metal2 s 312 34317 312 34317 4 wl0_86
port 977 nsew
rlabel metal2 s 312 29357 312 29357 4 wl1_74
port 954 nsew
rlabel metal2 s 312 28093 312 28093 4 wl0_71
port 947 nsew
rlabel metal2 s 312 37793 312 37793 4 wl1_95
port 996 nsew
rlabel metal2 s 312 38047 312 38047 4 wl1_96
port 998 nsew
rlabel metal2 s 312 27303 312 27303 4 wl0_69
port 943 nsew
rlabel metal2 s 312 37573 312 37573 4 wl0_95
port 995 nsew
rlabel metal2 s 312 30147 312 30147 4 wl1_76
port 958 nsew
rlabel metal2 s 312 35203 312 35203 4 wl0_89
port 983 nsew
rlabel metal2 s 312 34097 312 34097 4 wl1_86
port 978 nsew
rlabel metal2 s 312 32737 312 32737 4 wl0_82
port 969 nsew
rlabel metal2 s 312 37003 312 37003 4 wl1_93
port 992 nsew
rlabel metal2 s 312 30937 312 30937 4 wl1_78
port 962 nsew
rlabel metal2 s 312 29893 312 29893 4 wl1_75
port 956 nsew
rlabel metal2 s 312 28567 312 28567 4 wl1_72
port 950 nsew
rlabel metal2 s 312 27523 312 27523 4 wl1_69
port 944 nsew
rlabel metal2 s 312 33623 312 33623 4 wl0_85
port 975 nsew
rlabel metal2 s 312 29577 312 29577 4 wl0_74
port 953 nsew
rlabel metal2 s 312 33527 312 33527 4 wl0_84
port 973 nsew
rlabel metal2 s 312 34633 312 34633 4 wl1_87
port 980 nsew
rlabel metal2 s 312 34887 312 34887 4 wl1_88
port 982 nsew
rlabel metal2 s 312 26417 312 26417 4 wl0_66
port 937 nsew
rlabel metal2 s 312 15673 312 15673 4 wl1_39
port 884 nsew
rlabel metal2 s 312 24617 312 24617 4 wl1_62
port 930 nsew
rlabel metal2 s 312 15927 312 15927 4 wl1_40
port 886 nsew
rlabel metal2 s 312 20413 312 20413 4 wl1_51
port 908 nsew
rlabel metal2 s 312 19403 312 19403 4 wl0_49
port 903 nsew
rlabel metal2 s 312 19877 312 19877 4 wl1_50
port 906 nsew
rlabel metal2 s 312 25627 312 25627 4 wl0_64
port 933 nsew
rlabel metal2 s 312 17727 312 17727 4 wl0_44
port 893 nsew
rlabel metal2 s 312 16463 312 16463 4 wl1_41
port 888 nsew
rlabel metal2 s 312 25153 312 25153 4 wl1_63
port 932 nsew
rlabel metal2 s 312 18517 312 18517 4 wl0_46
port 897 nsew
rlabel metal2 s 312 22247 312 22247 4 wl1_56
port 918 nsew
rlabel metal2 s 312 25943 312 25943 4 wl1_65
port 936 nsew
rlabel metal2 s 312 24143 312 24143 4 wl0_61
port 927 nsew
rlabel metal2 s 312 22467 312 22467 4 wl0_56
port 917 nsew
rlabel metal2 s 312 18833 312 18833 4 wl1_47
port 900 nsew
rlabel metal2 s 312 24933 312 24933 4 wl0_63
port 931 nsew
rlabel metal2 s 312 21677 312 21677 4 wl0_54
port 913 nsew
rlabel metal2 s 312 14883 312 14883 4 wl1_37
port 880 nsew
rlabel metal2 s 312 16717 312 16717 4 wl1_42
port 890 nsew
rlabel metal2 s 312 23573 312 23573 4 wl1_59
port 924 nsew
rlabel metal2 s 312 21773 312 21773 4 wl0_55
port 915 nsew
rlabel metal2 s 312 23827 312 23827 4 wl1_60
port 926 nsew
rlabel metal2 s 312 17033 312 17033 4 wl0_43
port 891 nsew
rlabel metal2 s 312 16147 312 16147 4 wl0_40
port 885 nsew
rlabel metal2 s 312 23257 312 23257 4 wl0_58
port 921 nsew
rlabel metal2 s 312 25407 312 25407 4 wl1_64
port 934 nsew
rlabel metal2 s 312 17253 312 17253 4 wl1_43
port 892 nsew
rlabel metal2 s 312 20887 312 20887 4 wl0_52
port 909 nsew
rlabel metal2 s 312 18613 312 18613 4 wl0_47
port 899 nsew
rlabel metal2 s 312 16243 312 16243 4 wl0_41
port 887 nsew
rlabel metal2 s 312 17507 312 17507 4 wl1_44
port 894 nsew
rlabel metal2 s 312 13873 312 13873 4 wl0_35
port 875 nsew
rlabel metal2 s 312 20097 312 20097 4 wl0_50
port 905 nsew
rlabel metal2 s 312 15137 312 15137 4 wl1_38
port 882 nsew
rlabel metal2 s 312 14663 312 14663 4 wl0_37
port 879 nsew
rlabel metal2 s 312 15453 312 15453 4 wl0_39
port 883 nsew
rlabel metal2 s 312 19087 312 19087 4 wl1_48
port 902 nsew
rlabel metal2 s 312 15357 312 15357 4 wl0_38
port 881 nsew
rlabel metal2 s 312 19623 312 19623 4 wl1_49
port 904 nsew
rlabel metal2 s 312 19307 312 19307 4 wl0_48
port 901 nsew
rlabel metal2 s 312 21993 312 21993 4 wl1_55
port 916 nsew
rlabel metal2 s 312 23353 312 23353 4 wl0_59
port 923 nsew
rlabel metal2 s 312 23037 312 23037 4 wl1_58
port 922 nsew
rlabel metal2 s 312 22563 312 22563 4 wl0_57
port 919 nsew
rlabel metal2 s 312 14347 312 14347 4 wl1_36
port 878 nsew
rlabel metal2 s 312 13303 312 13303 4 wl1_33
port 872 nsew
rlabel metal2 s 312 21203 312 21203 4 wl1_53
port 912 nsew
rlabel metal2 s 312 17823 312 17823 4 wl0_45
port 895 nsew
rlabel metal2 s 312 13557 312 13557 4 wl1_34
port 874 nsew
rlabel metal2 s 312 21457 312 21457 4 wl1_54
port 914 nsew
rlabel metal2 s 312 18043 312 18043 4 wl1_45
port 896 nsew
rlabel metal2 s 312 25723 312 25723 4 wl0_65
port 935 nsew
rlabel metal2 s 312 18297 312 18297 4 wl1_46
port 898 nsew
rlabel metal2 s 312 24363 312 24363 4 wl1_61
port 928 nsew
rlabel metal2 s 312 16937 312 16937 4 wl0_42
port 889 nsew
rlabel metal2 s 312 22783 312 22783 4 wl1_57
port 920 nsew
rlabel metal2 s 312 14093 312 14093 4 wl1_35
port 876 nsew
rlabel metal2 s 312 14567 312 14567 4 wl0_36
port 877 nsew
rlabel metal2 s 312 20193 312 20193 4 wl0_51
port 907 nsew
rlabel metal2 s 312 24837 312 24837 4 wl0_62
port 929 nsew
rlabel metal2 s 312 20983 312 20983 4 wl0_53
port 911 nsew
rlabel metal2 s 312 24047 312 24047 4 wl0_60
port 925 nsew
rlabel metal2 s 312 13777 312 13777 4 wl0_34
port 873 nsew
rlabel metal2 s 312 20667 312 20667 4 wl1_52
port 910 nsew
rlabel metal2 s 312 1137 312 1137 4 wl0_2
port 809 nsew
rlabel metal2 s 312 3287 312 3287 4 wl1_8
port 822 nsew
rlabel metal2 s 312 1707 312 1707 4 wl1_4
port 814 nsew
rlabel metal2 s 312 4393 312 4393 4 wl0_11
port 827 nsew
rlabel metal2 s 312 2497 312 2497 4 wl1_6
port 818 nsew
rlabel metal2 s 312 9353 312 9353 4 wl1_23
port 852 nsew
rlabel metal2 s 312 6193 312 6193 4 wl1_15
port 836 nsew
rlabel metal2 s 312 9923 312 9923 4 wl0_25
port 855 nsew
rlabel metal2 s 312 1233 312 1233 4 wl0_3
port 811 nsew
rlabel metal2 s 312 9133 312 9133 4 wl0_23
port 851 nsew
rlabel metal2 s 312 5087 312 5087 4 wl0_12
port 829 nsew
rlabel metal2 s 312 10617 312 10617 4 wl0_26
port 857 nsew
rlabel metal2 s 312 7773 312 7773 4 wl1_19
port 844 nsew
rlabel metal2 s 312 6763 312 6763 4 wl0_17
port 839 nsew
rlabel metal2 s 312 917 312 917 4 wl1_2
port 810 nsew
rlabel metal2 s 312 5403 312 5403 4 wl1_13
port 832 nsew
rlabel metal2 s 312 1927 312 1927 4 wl0_4
port 813 nsew
rlabel metal2 s 312 10397 312 10397 4 wl1_26
port 858 nsew
rlabel metal2 s 312 7553 312 7553 4 wl0_19
port 843 nsew
rlabel metal2 s 312 11723 312 11723 4 wl1_29
port 864 nsew
rlabel metal2 s 312 4613 312 4613 4 wl1_11
port 828 nsew
rlabel metal2 s 312 12987 312 12987 4 wl0_32
port 869 nsew
rlabel metal2 s 312 6983 312 6983 4 wl1_17
port 840 nsew
rlabel metal2 s 312 6447 312 6447 4 wl1_16
port 838 nsew
rlabel metal2 s 312 3603 312 3603 4 wl0_9
port 823 nsew
rlabel metal2 s 312 12767 312 12767 4 wl1_32
port 870 nsew
rlabel metal2 s 312 2023 312 2023 4 wl0_5
port 815 nsew
rlabel metal2 s 312 11407 312 11407 4 wl0_28
port 861 nsew
rlabel metal2 s 312 8343 312 8343 4 wl0_21
port 847 nsew
rlabel metal2 s 312 3033 312 3033 4 wl1_7
port 820 nsew
rlabel metal2 s 312 10713 312 10713 4 wl0_27
port 859 nsew
rlabel metal2 s 312 8563 312 8563 4 wl1_21
port 848 nsew
rlabel metal2 s 312 11503 312 11503 4 wl0_29
port 863 nsew
rlabel metal2 s 312 8027 312 8027 4 wl1_20
port 846 nsew
rlabel metal2 s 312 10143 312 10143 4 wl1_25
port 856 nsew
rlabel metal2 s 312 5877 312 5877 4 wl0_14
port 833 nsew
rlabel metal2 s 312 2717 312 2717 4 wl0_6
port 817 nsew
rlabel metal2 s 312 10933 312 10933 4 wl1_27
port 860 nsew
rlabel metal2 s 312 2243 312 2243 4 wl1_5
port 816 nsew
rlabel metal2 s 312 11977 312 11977 4 wl1_30
port 866 nsew
rlabel metal2 s 312 4077 312 4077 4 wl1_10
port 826 nsew
rlabel metal2 s 312 12513 312 12513 4 wl1_31
port 868 nsew
rlabel metal2 s 312 13083 312 13083 4 wl0_33
port 871 nsew
rlabel metal2 s 312 7237 312 7237 4 wl1_18
port 842 nsew
rlabel metal2 s 312 2813 312 2813 4 wl0_7
port 819 nsew
rlabel metal2 s 312 5657 312 5657 4 wl1_14
port 834 nsew
rlabel metal2 s 312 9037 312 9037 4 wl0_22
port 849 nsew
rlabel metal2 s 312 11187 312 11187 4 wl1_28
port 862 nsew
rlabel metal2 s 312 3823 312 3823 4 wl1_9
port 824 nsew
rlabel metal2 s 312 663 312 663 4 wl1_1
port 808 nsew
rlabel metal2 s 312 3507 312 3507 4 wl0_8
port 821 nsew
rlabel metal2 s 312 8247 312 8247 4 wl0_20
port 845 nsew
rlabel metal2 s 312 6667 312 6667 4 wl0_16
port 837 nsew
rlabel metal2 s 312 4297 312 4297 4 wl0_10
port 825 nsew
rlabel metal2 s 312 12197 312 12197 4 wl0_30
port 865 nsew
rlabel metal2 s 312 4867 312 4867 4 wl1_12
port 830 nsew
rlabel metal2 s 312 443 312 443 4 wl0_1
port 807 nsew
rlabel metal2 s 312 5183 312 5183 4 wl0_13
port 831 nsew
rlabel metal2 s 312 9607 312 9607 4 wl1_24
port 854 nsew
rlabel metal2 s 312 7457 312 7457 4 wl0_18
port 841 nsew
rlabel metal2 s 312 5973 312 5973 4 wl0_15
port 835 nsew
rlabel metal2 s 312 1453 312 1453 4 wl1_3
port 812 nsew
rlabel metal2 s 312 8817 312 8817 4 wl1_22
port 850 nsew
rlabel metal2 s 312 12293 312 12293 4 wl0_31
port 867 nsew
rlabel metal2 s 312 9827 312 9827 4 wl0_24
port 853 nsew
rlabel metal2 s 384 7900 384 7900 4 gnd
port 2 nsew
rlabel metal2 s 384 8690 384 8690 4 gnd
port 2 nsew
rlabel metal2 s 384 18170 384 18170 4 gnd
port 2 nsew
rlabel metal2 s 384 22357 384 22357 4 gnd
port 2 nsew
rlabel metal2 s 384 20777 384 20777 4 gnd
port 2 nsew
rlabel metal2 s 384 19987 384 19987 4 gnd
port 2 nsew
rlabel metal2 s 384 2923 384 2923 4 gnd
port 2 nsew
rlabel metal2 s 384 7663 384 7663 4 gnd
port 2 nsew
rlabel metal2 s 384 18960 384 18960 4 gnd
port 2 nsew
rlabel metal2 s 384 9480 384 9480 4 gnd
port 2 nsew
rlabel metal2 s 384 11850 384 11850 4 gnd
port 2 nsew
rlabel metal2 s 384 16827 384 16827 4 gnd
port 2 nsew
rlabel metal2 s 384 22910 384 22910 4 gnd
port 2 nsew
rlabel metal2 s 384 11297 384 11297 4 gnd
port 2 nsew
rlabel metal2 s 384 13193 384 13193 4 gnd
port 2 nsew
rlabel metal2 s 384 21567 384 21567 4 gnd
port 2 nsew
rlabel metal2 s 384 2370 384 2370 4 gnd
port 2 nsew
rlabel metal2 s 384 16590 384 16590 4 gnd
port 2 nsew
rlabel metal2 s 384 26070 384 26070 4 gnd
port 2 nsew
rlabel metal2 s 384 5530 384 5530 4 gnd
port 2 nsew
rlabel metal2 s 384 13430 384 13430 4 gnd
port 2 nsew
rlabel metal2 s 384 25517 384 25517 4 gnd
port 2 nsew
rlabel metal2 s 384 1027 384 1027 4 gnd
port 2 nsew
rlabel metal2 s 384 8453 384 8453 4 gnd
port 2 nsew
rlabel metal2 s 384 9717 384 9717 4 gnd
port 2 nsew
rlabel metal2 s 384 23463 384 23463 4 gnd
port 2 nsew
rlabel metal2 s 384 14457 384 14457 4 gnd
port 2 nsew
rlabel metal2 s 384 7110 384 7110 4 gnd
port 2 nsew
rlabel metal2 s 384 21093 384 21093 4 gnd
port 2 nsew
rlabel metal2 s 384 22120 384 22120 4 gnd
port 2 nsew
rlabel metal2 s 384 21330 384 21330 4 gnd
port 2 nsew
rlabel metal2 s 384 3160 384 3160 4 gnd
port 2 nsew
rlabel metal2 s 384 3713 384 3713 4 gnd
port 2 nsew
rlabel metal2 s 384 25833 384 25833 4 gnd
port 2 nsew
rlabel metal2 s 384 10270 384 10270 4 gnd
port 2 nsew
rlabel metal2 s 384 15247 384 15247 4 gnd
port 2 nsew
rlabel metal2 s 384 553 384 553 4 gnd
port 2 nsew
rlabel metal2 s 384 11060 384 11060 4 gnd
port 2 nsew
rlabel metal2 s 384 23937 384 23937 4 gnd
port 2 nsew
rlabel metal2 s 384 17617 384 17617 4 gnd
port 2 nsew
rlabel metal2 s 384 8137 384 8137 4 gnd
port 2 nsew
rlabel metal2 s 384 15010 384 15010 4 gnd
port 2 nsew
rlabel metal2 s 384 15800 384 15800 4 gnd
port 2 nsew
rlabel metal2 s 384 18407 384 18407 4 gnd
port 2 nsew
rlabel metal2 s 384 17143 384 17143 4 gnd
port 2 nsew
rlabel metal2 s 384 25280 384 25280 4 gnd
port 2 nsew
rlabel metal2 s 384 4740 384 4740 4 gnd
port 2 nsew
rlabel metal2 s 384 9243 384 9243 4 gnd
port 2 nsew
rlabel metal2 s 384 5767 384 5767 4 gnd
port 2 nsew
rlabel metal2 s 384 7347 384 7347 4 gnd
port 2 nsew
rlabel metal2 s 384 19750 384 19750 4 gnd
port 2 nsew
rlabel metal2 s 384 12640 384 12640 4 gnd
port 2 nsew
rlabel metal2 s 384 24253 384 24253 4 gnd
port 2 nsew
rlabel metal2 s 384 4503 384 4503 4 gnd
port 2 nsew
rlabel metal2 s 384 22673 384 22673 4 gnd
port 2 nsew
rlabel metal2 s 384 6320 384 6320 4 gnd
port 2 nsew
rlabel metal2 s 384 18723 384 18723 4 gnd
port 2 nsew
rlabel metal2 s 384 21883 384 21883 4 gnd
port 2 nsew
rlabel metal2 s 384 4187 384 4187 4 gnd
port 2 nsew
rlabel metal2 s 384 14220 384 14220 4 gnd
port 2 nsew
rlabel metal2 s 384 10507 384 10507 4 gnd
port 2 nsew
rlabel metal2 s 384 11613 384 11613 4 gnd
port 2 nsew
rlabel metal2 s 384 8927 384 8927 4 gnd
port 2 nsew
rlabel metal2 s 384 6873 384 6873 4 gnd
port 2 nsew
rlabel metal2 s 384 2607 384 2607 4 gnd
port 2 nsew
rlabel metal2 s 384 1580 384 1580 4 gnd
port 2 nsew
rlabel metal2 s 384 17933 384 17933 4 gnd
port 2 nsew
rlabel metal2 s 384 19197 384 19197 4 gnd
port 2 nsew
rlabel metal2 s 384 12403 384 12403 4 gnd
port 2 nsew
rlabel metal2 s 384 1343 384 1343 4 gnd
port 2 nsew
rlabel metal2 s 384 15563 384 15563 4 gnd
port 2 nsew
rlabel metal2 s 384 20540 384 20540 4 gnd
port 2 nsew
rlabel metal2 s 384 6083 384 6083 4 gnd
port 2 nsew
rlabel metal2 s 384 4977 384 4977 4 gnd
port 2 nsew
rlabel metal2 s 384 17380 384 17380 4 gnd
port 2 nsew
rlabel metal2 s 384 12087 384 12087 4 gnd
port 2 nsew
rlabel metal2 s 384 790 384 790 4 gnd
port 2 nsew
rlabel metal2 s 384 23700 384 23700 4 gnd
port 2 nsew
rlabel metal2 s 384 25043 384 25043 4 gnd
port 2 nsew
rlabel metal2 s 384 2133 384 2133 4 gnd
port 2 nsew
rlabel metal2 s 384 1817 384 1817 4 gnd
port 2 nsew
rlabel metal2 s 384 3397 384 3397 4 gnd
port 2 nsew
rlabel metal2 s 384 13983 384 13983 4 gnd
port 2 nsew
rlabel metal2 s 384 5293 384 5293 4 gnd
port 2 nsew
rlabel metal2 s 384 6557 384 6557 4 gnd
port 2 nsew
rlabel metal2 s 384 24727 384 24727 4 gnd
port 2 nsew
rlabel metal2 s 384 10033 384 10033 4 gnd
port 2 nsew
rlabel metal2 s 384 10823 384 10823 4 gnd
port 2 nsew
rlabel metal2 s 384 3950 384 3950 4 gnd
port 2 nsew
rlabel metal2 s 384 13667 384 13667 4 gnd
port 2 nsew
rlabel metal2 s 384 14773 384 14773 4 gnd
port 2 nsew
rlabel metal2 s 384 20303 384 20303 4 gnd
port 2 nsew
rlabel metal2 s 384 24490 384 24490 4 gnd
port 2 nsew
rlabel metal2 s 384 23147 384 23147 4 gnd
port 2 nsew
rlabel metal2 s 384 16037 384 16037 4 gnd
port 2 nsew
rlabel metal2 s 384 16353 384 16353 4 gnd
port 2 nsew
rlabel metal2 s 384 19513 384 19513 4 gnd
port 2 nsew
rlabel metal2 s 384 12877 384 12877 4 gnd
port 2 nsew
rlabel metal3 s 312 229 312 229 4 vdd
port 1 nsew
rlabel metal3 s 312 51911 312 51911 4 vdd
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 624 52140
string GDS_END 4319350
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 4235318
<< end >>
