magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< pwell >>
rect -10 -26 76 1246
rect 266 564 287 613
rect 494 -26 580 1246
<< locali >>
rect 16 0 50 1220
rect 520 0 554 1220
<< metal1 >>
rect 16 1213 554 1220
rect 16 1161 59 1213
rect 111 1161 139 1213
rect 191 1161 219 1213
rect 271 1161 299 1213
rect 351 1161 379 1213
rect 431 1161 459 1213
rect 511 1161 554 1213
rect 16 1154 554 1161
rect 16 126 50 1154
rect 78 66 114 1094
rect 142 126 176 1154
rect 204 66 240 1094
rect 268 126 302 1154
rect 330 66 366 1094
rect 394 126 428 1154
rect 456 66 492 1094
rect 520 126 554 1154
rect 66 59 504 66
rect 66 7 99 59
rect 151 7 179 59
rect 231 7 259 59
rect 311 7 339 59
rect 391 7 419 59
rect 471 7 504 59
rect 66 0 504 7
<< via1 >>
rect 59 1161 111 1213
rect 139 1161 191 1213
rect 219 1161 271 1213
rect 299 1161 351 1213
rect 379 1161 431 1213
rect 459 1161 511 1213
rect 99 7 151 59
rect 179 7 231 59
rect 259 7 311 59
rect 339 7 391 59
rect 419 7 471 59
<< metal2 >>
rect 16 1215 554 1220
rect 16 1159 57 1215
rect 113 1159 137 1215
rect 193 1159 217 1215
rect 273 1159 297 1215
rect 353 1159 377 1215
rect 433 1159 457 1215
rect 513 1159 554 1215
rect 16 1154 554 1159
rect 16 126 50 1154
rect 78 66 114 1094
rect 142 126 176 1154
rect 204 66 240 1094
rect 268 126 302 1154
rect 330 66 366 1094
rect 394 126 428 1154
rect 456 66 492 1094
rect 520 126 554 1154
rect 66 61 504 66
rect 66 5 97 61
rect 153 5 177 61
rect 233 5 257 61
rect 313 5 337 61
rect 393 5 417 61
rect 473 5 504 61
rect 66 0 504 5
<< via2 >>
rect 57 1213 113 1215
rect 57 1161 59 1213
rect 59 1161 111 1213
rect 111 1161 113 1213
rect 57 1159 113 1161
rect 137 1213 193 1215
rect 137 1161 139 1213
rect 139 1161 191 1213
rect 191 1161 193 1213
rect 137 1159 193 1161
rect 217 1213 273 1215
rect 217 1161 219 1213
rect 219 1161 271 1213
rect 271 1161 273 1213
rect 217 1159 273 1161
rect 297 1213 353 1215
rect 297 1161 299 1213
rect 299 1161 351 1213
rect 351 1161 353 1213
rect 297 1159 353 1161
rect 377 1213 433 1215
rect 377 1161 379 1213
rect 379 1161 431 1213
rect 431 1161 433 1213
rect 377 1159 433 1161
rect 457 1213 513 1215
rect 457 1161 459 1213
rect 459 1161 511 1213
rect 511 1161 513 1213
rect 457 1159 513 1161
rect 97 59 153 61
rect 97 7 99 59
rect 99 7 151 59
rect 151 7 153 59
rect 97 5 153 7
rect 177 59 233 61
rect 177 7 179 59
rect 179 7 231 59
rect 231 7 233 59
rect 177 5 233 7
rect 257 59 313 61
rect 257 7 259 59
rect 259 7 311 59
rect 311 7 313 59
rect 257 5 313 7
rect 337 59 393 61
rect 337 7 339 59
rect 339 7 391 59
rect 391 7 393 59
rect 337 5 393 7
rect 417 59 473 61
rect 417 7 419 59
rect 419 7 471 59
rect 471 7 473 59
rect 417 5 473 7
<< metal3 >>
rect 0 1215 570 1220
rect 0 1159 57 1215
rect 113 1159 137 1215
rect 193 1159 217 1215
rect 273 1159 297 1215
rect 353 1159 377 1215
rect 433 1159 457 1215
rect 513 1159 570 1215
rect 0 1154 570 1159
rect 0 1141 66 1154
rect 0 1077 1 1141
rect 65 1077 66 1141
rect 252 1141 318 1154
rect 0 1015 66 1077
rect 0 951 1 1015
rect 65 951 66 1015
rect 0 889 66 951
rect 0 825 1 889
rect 65 825 66 889
rect 0 763 66 825
rect 0 699 1 763
rect 65 699 66 763
rect 0 637 66 699
rect 0 573 1 637
rect 65 573 66 637
rect 0 511 66 573
rect 0 447 1 511
rect 65 447 66 511
rect 0 385 66 447
rect 0 321 1 385
rect 65 321 66 385
rect 0 259 66 321
rect 0 195 1 259
rect 65 195 66 259
rect 0 126 66 195
rect 126 1078 192 1094
rect 126 1014 127 1078
rect 191 1014 192 1078
rect 126 952 192 1014
rect 126 888 127 952
rect 191 888 192 952
rect 126 826 192 888
rect 126 762 127 826
rect 191 762 192 826
rect 126 700 192 762
rect 126 636 127 700
rect 191 636 192 700
rect 126 574 192 636
rect 126 510 127 574
rect 191 510 192 574
rect 126 448 192 510
rect 126 384 127 448
rect 191 384 192 448
rect 126 322 192 384
rect 126 258 127 322
rect 191 258 192 322
rect 126 196 192 258
rect 126 132 127 196
rect 191 132 192 196
rect 126 66 192 132
rect 252 1077 253 1141
rect 317 1077 318 1141
rect 504 1141 570 1154
rect 252 1015 318 1077
rect 252 951 253 1015
rect 317 951 318 1015
rect 252 889 318 951
rect 252 825 253 889
rect 317 825 318 889
rect 252 763 318 825
rect 252 699 253 763
rect 317 699 318 763
rect 252 637 318 699
rect 252 573 253 637
rect 317 573 318 637
rect 252 511 318 573
rect 252 447 253 511
rect 317 447 318 511
rect 252 385 318 447
rect 252 321 253 385
rect 317 321 318 385
rect 252 259 318 321
rect 252 195 253 259
rect 317 195 318 259
rect 252 126 318 195
rect 378 1078 444 1094
rect 378 1014 379 1078
rect 443 1014 444 1078
rect 378 952 444 1014
rect 378 888 379 952
rect 443 888 444 952
rect 378 826 444 888
rect 378 762 379 826
rect 443 762 444 826
rect 378 700 444 762
rect 378 636 379 700
rect 443 636 444 700
rect 378 574 444 636
rect 378 510 379 574
rect 443 510 444 574
rect 378 448 444 510
rect 378 384 379 448
rect 443 384 444 448
rect 378 322 444 384
rect 378 258 379 322
rect 443 258 444 322
rect 378 196 444 258
rect 378 132 379 196
rect 443 132 444 196
rect 378 66 444 132
rect 504 1077 505 1141
rect 569 1077 570 1141
rect 504 1015 570 1077
rect 504 951 505 1015
rect 569 951 570 1015
rect 504 889 570 951
rect 504 825 505 889
rect 569 825 570 889
rect 504 763 570 825
rect 504 699 505 763
rect 569 699 570 763
rect 504 637 570 699
rect 504 573 505 637
rect 569 573 570 637
rect 504 511 570 573
rect 504 447 505 511
rect 569 447 570 511
rect 504 385 570 447
rect 504 321 505 385
rect 569 321 570 385
rect 504 259 570 321
rect 504 195 505 259
rect 569 195 570 259
rect 504 126 570 195
rect 66 61 504 66
rect 66 5 97 61
rect 153 5 177 61
rect 233 5 257 61
rect 313 5 337 61
rect 393 5 417 61
rect 473 5 504 61
rect 66 0 504 5
<< via3 >>
rect 1 1077 65 1141
rect 1 951 65 1015
rect 1 825 65 889
rect 1 699 65 763
rect 1 573 65 637
rect 1 447 65 511
rect 1 321 65 385
rect 1 195 65 259
rect 127 1014 191 1078
rect 127 888 191 952
rect 127 762 191 826
rect 127 636 191 700
rect 127 510 191 574
rect 127 384 191 448
rect 127 258 191 322
rect 127 132 191 196
rect 253 1077 317 1141
rect 253 951 317 1015
rect 253 825 317 889
rect 253 699 317 763
rect 253 573 317 637
rect 253 447 317 511
rect 253 321 317 385
rect 253 195 317 259
rect 379 1014 443 1078
rect 379 888 443 952
rect 379 762 443 826
rect 379 636 443 700
rect 379 510 443 574
rect 379 384 443 448
rect 379 258 443 322
rect 379 132 443 196
rect 505 1077 569 1141
rect 505 951 569 1015
rect 505 825 569 889
rect 505 699 569 763
rect 505 573 569 637
rect 505 447 569 511
rect 505 321 569 385
rect 505 195 569 259
<< metal4 >>
rect 0 1141 66 1220
rect 0 1077 1 1141
rect 65 1077 66 1141
rect 0 1015 66 1077
rect 0 951 1 1015
rect 65 951 66 1015
rect 0 889 66 951
rect 0 825 1 889
rect 65 825 66 889
rect 0 763 66 825
rect 0 699 1 763
rect 65 699 66 763
rect 0 637 66 699
rect 0 573 1 637
rect 65 573 66 637
rect 0 511 66 573
rect 0 447 1 511
rect 65 447 66 511
rect 0 385 66 447
rect 0 321 1 385
rect 65 321 66 385
rect 0 259 66 321
rect 0 195 1 259
rect 65 195 66 259
rect 0 66 66 195
rect 126 1078 192 1154
rect 126 1014 127 1078
rect 191 1014 192 1078
rect 126 952 192 1014
rect 126 888 127 952
rect 191 888 192 952
rect 126 826 192 888
rect 126 762 127 826
rect 191 762 192 826
rect 126 700 192 762
rect 126 636 127 700
rect 191 636 192 700
rect 126 574 192 636
rect 126 510 127 574
rect 191 510 192 574
rect 126 448 192 510
rect 126 384 127 448
rect 191 384 192 448
rect 126 322 192 384
rect 126 258 127 322
rect 191 258 192 322
rect 126 196 192 258
rect 126 132 127 196
rect 191 132 192 196
rect 126 0 192 132
rect 252 1141 318 1220
rect 252 1077 253 1141
rect 317 1077 318 1141
rect 252 1015 318 1077
rect 252 951 253 1015
rect 317 951 318 1015
rect 252 889 318 951
rect 252 825 253 889
rect 317 825 318 889
rect 252 763 318 825
rect 252 699 253 763
rect 317 699 318 763
rect 252 637 318 699
rect 252 573 253 637
rect 317 573 318 637
rect 252 511 318 573
rect 252 447 253 511
rect 317 447 318 511
rect 252 385 318 447
rect 252 321 253 385
rect 317 321 318 385
rect 252 259 318 321
rect 252 195 253 259
rect 317 195 318 259
rect 252 66 318 195
rect 378 1078 444 1154
rect 378 1014 379 1078
rect 443 1014 444 1078
rect 378 952 444 1014
rect 378 888 379 952
rect 443 888 444 952
rect 378 826 444 888
rect 378 762 379 826
rect 443 762 444 826
rect 378 700 444 762
rect 378 636 379 700
rect 443 636 444 700
rect 378 574 444 636
rect 378 510 379 574
rect 443 510 444 574
rect 378 448 444 510
rect 378 384 379 448
rect 443 384 444 448
rect 378 322 444 384
rect 378 258 379 322
rect 443 258 444 322
rect 378 196 444 258
rect 378 132 379 196
rect 443 132 444 196
rect 378 0 444 132
rect 504 1141 570 1220
rect 504 1077 505 1141
rect 569 1077 570 1141
rect 504 1015 570 1077
rect 504 951 505 1015
rect 569 951 570 1015
rect 504 889 570 951
rect 504 825 505 889
rect 569 825 570 889
rect 504 763 570 825
rect 504 699 505 763
rect 569 699 570 763
rect 504 637 570 699
rect 504 573 505 637
rect 569 573 570 637
rect 504 511 570 573
rect 504 447 505 511
rect 569 447 570 511
rect 504 385 570 447
rect 504 321 505 385
rect 569 321 570 385
rect 504 259 570 321
rect 504 195 505 259
rect 569 195 570 259
rect 504 66 570 195
<< labels >>
flabel metal2 s 149 262 168 282 0 FreeSans 200 0 0 0 C0
port 1 nsew
flabel metal2 s 330 72 366 108 0 FreeSans 200 0 0 0 C1
port 2 nsew
flabel pwell s 266 564 287 613 0 FreeSans 400 0 0 0 SUB
port 3 nsew
<< properties >>
string GDS_END 55600
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 46816
string path 1.650 0.825 12.600 0.825 
string device primitive
<< end >>
