magic
tech sky130B
timestamp 1683767628
<< properties >>
string GDS_END 15506366
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 15503610
<< end >>
