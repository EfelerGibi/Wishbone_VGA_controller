magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< locali >>
rect 243 961 559 980
rect 243 927 255 961
rect 289 927 337 961
rect 371 927 431 961
rect 465 927 513 961
rect 547 927 559 961
rect 243 889 559 927
rect 120 823 186 889
rect 243 855 255 889
rect 289 855 337 889
rect 371 855 431 889
rect 465 855 513 889
rect 547 855 559 889
rect 243 841 559 855
rect 616 823 682 889
rect 120 795 160 823
rect 642 795 682 823
rect 41 759 160 795
rect 41 725 60 759
rect 94 725 160 759
rect 41 687 160 725
rect 41 653 60 687
rect 94 653 160 687
rect 41 615 160 653
rect 41 581 60 615
rect 94 581 160 615
rect 41 543 160 581
rect 41 509 60 543
rect 94 509 160 543
rect 41 471 160 509
rect 41 437 60 471
rect 94 437 160 471
rect 41 399 160 437
rect 41 365 60 399
rect 94 365 160 399
rect 41 327 160 365
rect 41 293 60 327
rect 94 293 160 327
rect 41 255 160 293
rect 41 221 60 255
rect 94 221 160 255
rect 41 185 160 221
rect 642 759 761 795
rect 642 725 708 759
rect 742 725 761 759
rect 642 687 761 725
rect 642 653 708 687
rect 742 653 761 687
rect 642 615 761 653
rect 642 581 708 615
rect 742 581 761 615
rect 642 543 761 581
rect 642 509 708 543
rect 742 509 761 543
rect 642 471 761 509
rect 642 437 708 471
rect 742 437 761 471
rect 642 399 761 437
rect 642 365 708 399
rect 742 365 761 399
rect 642 327 761 365
rect 642 293 708 327
rect 742 293 761 327
rect 642 255 761 293
rect 642 221 708 255
rect 742 221 761 255
rect 642 185 761 221
rect 120 157 160 185
rect 642 157 682 185
rect 120 91 186 157
rect 243 125 559 139
rect 243 91 255 125
rect 289 91 337 125
rect 371 91 431 125
rect 465 91 513 125
rect 547 91 559 125
rect 616 91 682 157
rect 243 53 559 91
rect 243 19 255 53
rect 289 19 337 53
rect 371 19 431 53
rect 465 19 513 53
rect 547 19 559 53
rect 243 0 559 19
<< viali >>
rect 255 927 289 961
rect 337 927 371 961
rect 431 927 465 961
rect 513 927 547 961
rect 255 855 289 889
rect 337 855 371 889
rect 431 855 465 889
rect 513 855 547 889
rect 60 725 94 759
rect 60 653 94 687
rect 60 581 94 615
rect 60 509 94 543
rect 60 437 94 471
rect 60 365 94 399
rect 60 293 94 327
rect 60 221 94 255
rect 708 725 742 759
rect 708 653 742 687
rect 708 581 742 615
rect 708 509 742 543
rect 708 437 742 471
rect 708 365 742 399
rect 708 293 742 327
rect 708 221 742 255
rect 255 91 289 125
rect 337 91 371 125
rect 431 91 465 125
rect 513 91 547 125
rect 255 19 289 53
rect 337 19 371 53
rect 431 19 465 53
rect 513 19 547 53
<< obsli1 >>
rect 212 185 246 795
rect 298 185 332 795
rect 384 185 418 795
rect 470 185 504 795
rect 556 185 590 795
<< metal1 >>
rect 243 961 559 980
rect 243 927 255 961
rect 289 927 337 961
rect 371 927 431 961
rect 465 927 513 961
rect 547 927 559 961
rect 243 889 559 927
rect 243 855 255 889
rect 289 855 337 889
rect 371 855 431 889
rect 465 855 513 889
rect 547 855 559 889
rect 243 843 559 855
rect 41 759 100 771
rect 41 725 60 759
rect 94 725 100 759
rect 41 687 100 725
rect 41 653 60 687
rect 94 653 100 687
rect 41 615 100 653
rect 41 581 60 615
rect 94 581 100 615
rect 41 543 100 581
rect 41 509 60 543
rect 94 509 100 543
rect 41 471 100 509
rect 41 437 60 471
rect 94 437 100 471
rect 41 399 100 437
rect 41 365 60 399
rect 94 365 100 399
rect 41 327 100 365
rect 41 293 60 327
rect 94 293 100 327
rect 41 255 100 293
rect 41 221 60 255
rect 94 221 100 255
rect 41 209 100 221
rect 702 759 761 771
rect 702 725 708 759
rect 742 725 761 759
rect 702 687 761 725
rect 702 653 708 687
rect 742 653 761 687
rect 702 615 761 653
rect 702 581 708 615
rect 742 581 761 615
rect 702 543 761 581
rect 702 509 708 543
rect 742 509 761 543
rect 702 471 761 509
rect 702 437 708 471
rect 742 437 761 471
rect 702 399 761 437
rect 702 365 708 399
rect 742 365 761 399
rect 702 327 761 365
rect 702 293 708 327
rect 742 293 761 327
rect 702 255 761 293
rect 702 221 708 255
rect 742 221 761 255
rect 702 209 761 221
rect 243 125 559 137
rect 243 91 255 125
rect 289 91 337 125
rect 371 91 431 125
rect 465 91 513 125
rect 547 91 559 125
rect 243 53 559 91
rect 243 19 255 53
rect 289 19 337 53
rect 371 19 431 53
rect 465 19 513 53
rect 547 19 559 53
rect 243 0 559 19
<< obsm1 >>
rect 203 209 255 771
rect 289 209 341 771
rect 375 209 427 771
rect 461 209 513 771
rect 547 209 599 771
<< metal2 >>
rect 14 515 788 771
rect 14 209 788 465
<< labels >>
rlabel viali s 708 725 742 759 6 BULK
port 4 nsew
rlabel viali s 708 653 742 687 6 BULK
port 4 nsew
rlabel viali s 708 581 742 615 6 BULK
port 4 nsew
rlabel viali s 708 509 742 543 6 BULK
port 4 nsew
rlabel viali s 708 437 742 471 6 BULK
port 4 nsew
rlabel viali s 708 365 742 399 6 BULK
port 4 nsew
rlabel viali s 708 293 742 327 6 BULK
port 4 nsew
rlabel viali s 708 221 742 255 6 BULK
port 4 nsew
rlabel viali s 60 725 94 759 6 BULK
port 4 nsew
rlabel viali s 60 653 94 687 6 BULK
port 4 nsew
rlabel viali s 60 581 94 615 6 BULK
port 4 nsew
rlabel viali s 60 509 94 543 6 BULK
port 4 nsew
rlabel viali s 60 437 94 471 6 BULK
port 4 nsew
rlabel viali s 60 365 94 399 6 BULK
port 4 nsew
rlabel viali s 60 293 94 327 6 BULK
port 4 nsew
rlabel viali s 60 221 94 255 6 BULK
port 4 nsew
rlabel locali s 642 795 682 823 6 BULK
port 4 nsew
rlabel locali s 642 185 761 795 6 BULK
port 4 nsew
rlabel locali s 642 157 682 185 6 BULK
port 4 nsew
rlabel locali s 616 823 682 889 6 BULK
port 4 nsew
rlabel locali s 616 91 682 157 6 BULK
port 4 nsew
rlabel locali s 120 823 186 889 6 BULK
port 4 nsew
rlabel locali s 120 795 160 823 6 BULK
port 4 nsew
rlabel locali s 120 157 160 185 6 BULK
port 4 nsew
rlabel locali s 120 91 186 157 6 BULK
port 4 nsew
rlabel locali s 41 185 160 795 6 BULK
port 4 nsew
rlabel metal1 s 702 209 761 771 6 BULK
port 4 nsew
rlabel metal1 s 41 209 100 771 6 BULK
port 4 nsew
rlabel metal2 s 14 515 788 771 6 DRAIN
port 1 nsew
rlabel viali s 513 927 547 961 6 GATE
port 2 nsew
rlabel viali s 513 855 547 889 6 GATE
port 2 nsew
rlabel viali s 513 91 547 125 6 GATE
port 2 nsew
rlabel viali s 513 19 547 53 6 GATE
port 2 nsew
rlabel viali s 431 927 465 961 6 GATE
port 2 nsew
rlabel viali s 431 855 465 889 6 GATE
port 2 nsew
rlabel viali s 431 91 465 125 6 GATE
port 2 nsew
rlabel viali s 431 19 465 53 6 GATE
port 2 nsew
rlabel viali s 337 927 371 961 6 GATE
port 2 nsew
rlabel viali s 337 855 371 889 6 GATE
port 2 nsew
rlabel viali s 337 91 371 125 6 GATE
port 2 nsew
rlabel viali s 337 19 371 53 6 GATE
port 2 nsew
rlabel viali s 255 927 289 961 6 GATE
port 2 nsew
rlabel viali s 255 855 289 889 6 GATE
port 2 nsew
rlabel viali s 255 91 289 125 6 GATE
port 2 nsew
rlabel viali s 255 19 289 53 6 GATE
port 2 nsew
rlabel locali s 243 841 559 980 6 GATE
port 2 nsew
rlabel locali s 243 0 559 139 6 GATE
port 2 nsew
rlabel metal1 s 243 843 559 980 6 GATE
port 2 nsew
rlabel metal1 s 243 0 559 137 6 GATE
port 2 nsew
rlabel metal2 s 14 209 788 465 6 SOURCE
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 802 980
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9754396
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9734030
string device primitive
<< end >>