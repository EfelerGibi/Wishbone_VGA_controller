magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 1 21 1115 203
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 167 47 197 177
rect 251 47 281 177
rect 335 47 365 177
rect 419 47 449 177
rect 503 47 533 177
rect 587 47 617 177
rect 671 47 701 177
rect 755 47 785 177
rect 839 47 869 177
rect 923 47 953 177
rect 1007 47 1037 177
<< scpmoshvt >>
rect 83 297 113 497
rect 167 297 197 497
rect 251 297 281 497
rect 335 297 365 497
rect 419 297 449 497
rect 503 297 533 497
rect 587 297 617 497
rect 671 297 701 497
rect 755 297 785 497
rect 839 297 869 497
rect 923 297 953 497
rect 1007 297 1037 497
<< ndiff >>
rect 27 163 83 177
rect 27 129 39 163
rect 73 129 83 163
rect 27 95 83 129
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 167 177
rect 113 129 123 163
rect 157 129 167 163
rect 113 95 167 129
rect 113 61 123 95
rect 157 61 167 95
rect 113 47 167 61
rect 197 95 251 177
rect 197 61 207 95
rect 241 61 251 95
rect 197 47 251 61
rect 281 163 335 177
rect 281 129 291 163
rect 325 129 335 163
rect 281 95 335 129
rect 281 61 291 95
rect 325 61 335 95
rect 281 47 335 61
rect 365 95 419 177
rect 365 61 375 95
rect 409 61 419 95
rect 365 47 419 61
rect 449 163 503 177
rect 449 129 459 163
rect 493 129 503 163
rect 449 95 503 129
rect 449 61 459 95
rect 493 61 503 95
rect 449 47 503 61
rect 533 95 587 177
rect 533 61 543 95
rect 577 61 587 95
rect 533 47 587 61
rect 617 163 671 177
rect 617 129 627 163
rect 661 129 671 163
rect 617 95 671 129
rect 617 61 627 95
rect 661 61 671 95
rect 617 47 671 61
rect 701 95 755 177
rect 701 61 711 95
rect 745 61 755 95
rect 701 47 755 61
rect 785 163 839 177
rect 785 129 795 163
rect 829 129 839 163
rect 785 95 839 129
rect 785 61 795 95
rect 829 61 839 95
rect 785 47 839 61
rect 869 95 923 177
rect 869 61 879 95
rect 913 61 923 95
rect 869 47 923 61
rect 953 163 1007 177
rect 953 129 963 163
rect 997 129 1007 163
rect 953 95 1007 129
rect 953 61 963 95
rect 997 61 1007 95
rect 953 47 1007 61
rect 1037 95 1089 177
rect 1037 61 1047 95
rect 1081 61 1089 95
rect 1037 47 1089 61
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 341 83 375
rect 27 307 39 341
rect 73 307 83 341
rect 27 297 83 307
rect 113 477 167 497
rect 113 443 123 477
rect 157 443 167 477
rect 113 409 167 443
rect 113 375 123 409
rect 157 375 167 409
rect 113 297 167 375
rect 197 477 251 497
rect 197 443 207 477
rect 241 443 251 477
rect 197 409 251 443
rect 197 375 207 409
rect 241 375 251 409
rect 197 341 251 375
rect 197 307 207 341
rect 241 307 251 341
rect 197 297 251 307
rect 281 477 335 497
rect 281 443 291 477
rect 325 443 335 477
rect 281 409 335 443
rect 281 375 291 409
rect 325 375 335 409
rect 281 297 335 375
rect 365 477 419 497
rect 365 443 375 477
rect 409 443 419 477
rect 365 409 419 443
rect 365 375 375 409
rect 409 375 419 409
rect 365 341 419 375
rect 365 307 375 341
rect 409 307 419 341
rect 365 297 419 307
rect 449 341 503 497
rect 449 307 459 341
rect 493 307 503 341
rect 449 297 503 307
rect 533 477 587 497
rect 533 443 543 477
rect 577 443 587 477
rect 533 409 587 443
rect 533 375 543 409
rect 577 375 587 409
rect 533 297 587 375
rect 617 477 671 497
rect 617 443 627 477
rect 661 443 671 477
rect 617 409 671 443
rect 617 375 627 409
rect 661 375 671 409
rect 617 341 671 375
rect 617 307 627 341
rect 661 307 671 341
rect 617 297 671 307
rect 701 409 755 497
rect 701 375 711 409
rect 745 375 755 409
rect 701 297 755 375
rect 785 477 839 497
rect 785 443 795 477
rect 829 443 839 477
rect 785 297 839 443
rect 869 409 923 497
rect 869 375 879 409
rect 913 375 923 409
rect 869 297 923 375
rect 953 477 1007 497
rect 953 443 963 477
rect 997 443 1007 477
rect 953 297 1007 443
rect 1037 477 1089 497
rect 1037 443 1047 477
rect 1081 443 1089 477
rect 1037 297 1089 443
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 123 129 157 163
rect 123 61 157 95
rect 207 61 241 95
rect 291 129 325 163
rect 291 61 325 95
rect 375 61 409 95
rect 459 129 493 163
rect 459 61 493 95
rect 543 61 577 95
rect 627 129 661 163
rect 627 61 661 95
rect 711 61 745 95
rect 795 129 829 163
rect 795 61 829 95
rect 879 61 913 95
rect 963 129 997 163
rect 963 61 997 95
rect 1047 61 1081 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 123 443 157 477
rect 123 375 157 409
rect 207 443 241 477
rect 207 375 241 409
rect 207 307 241 341
rect 291 443 325 477
rect 291 375 325 409
rect 375 443 409 477
rect 375 375 409 409
rect 375 307 409 341
rect 459 307 493 341
rect 543 443 577 477
rect 543 375 577 409
rect 627 443 661 477
rect 627 375 661 409
rect 627 307 661 341
rect 711 375 745 409
rect 795 443 829 477
rect 879 375 913 409
rect 963 443 997 477
rect 1047 443 1081 477
<< poly >>
rect 83 497 113 523
rect 167 497 197 523
rect 251 497 281 523
rect 335 497 365 523
rect 419 497 449 523
rect 503 497 533 523
rect 587 497 617 523
rect 671 497 701 523
rect 755 497 785 523
rect 839 497 869 523
rect 923 497 953 523
rect 1007 497 1037 523
rect 83 265 113 297
rect 167 265 197 297
rect 251 265 281 297
rect 335 265 365 297
rect 83 249 365 265
rect 83 215 99 249
rect 133 215 167 249
rect 201 215 235 249
rect 269 215 303 249
rect 337 215 365 249
rect 83 199 365 215
rect 83 177 113 199
rect 167 177 197 199
rect 251 177 281 199
rect 335 177 365 199
rect 419 265 449 297
rect 503 265 533 297
rect 587 265 617 297
rect 419 249 617 265
rect 419 215 435 249
rect 469 215 503 249
rect 537 215 617 249
rect 419 199 617 215
rect 419 177 449 199
rect 503 177 533 199
rect 587 177 617 199
rect 671 265 701 297
rect 755 265 785 297
rect 839 265 869 297
rect 923 265 953 297
rect 1007 265 1037 297
rect 671 249 953 265
rect 671 215 823 249
rect 857 215 891 249
rect 925 215 953 249
rect 671 199 953 215
rect 999 249 1065 265
rect 999 215 1015 249
rect 1049 215 1065 249
rect 999 199 1065 215
rect 671 177 701 199
rect 755 177 785 199
rect 839 177 869 199
rect 923 177 953 199
rect 1007 177 1037 199
rect 83 21 113 47
rect 167 21 197 47
rect 251 21 281 47
rect 335 21 365 47
rect 419 21 449 47
rect 503 21 533 47
rect 587 21 617 47
rect 671 21 701 47
rect 755 21 785 47
rect 839 21 869 47
rect 923 21 953 47
rect 1007 21 1037 47
<< polycont >>
rect 99 215 133 249
rect 167 215 201 249
rect 235 215 269 249
rect 303 215 337 249
rect 435 215 469 249
rect 503 215 537 249
rect 823 215 857 249
rect 891 215 925 249
rect 1015 215 1049 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 30 477 81 493
rect 30 443 39 477
rect 73 443 81 477
rect 30 409 81 443
rect 30 375 39 409
rect 73 375 81 409
rect 30 341 81 375
rect 115 477 165 527
rect 115 443 123 477
rect 157 443 165 477
rect 115 409 165 443
rect 115 375 123 409
rect 157 375 165 409
rect 115 359 165 375
rect 199 477 249 493
rect 199 443 207 477
rect 241 443 249 477
rect 199 409 249 443
rect 199 375 207 409
rect 241 375 249 409
rect 30 307 39 341
rect 73 325 81 341
rect 199 341 249 375
rect 283 477 333 527
rect 283 443 291 477
rect 325 443 333 477
rect 283 409 333 443
rect 283 375 291 409
rect 325 375 333 409
rect 283 359 333 375
rect 367 477 585 493
rect 367 443 375 477
rect 409 459 543 477
rect 409 443 489 459
rect 367 425 489 443
rect 523 443 543 459
rect 577 443 585 477
rect 523 425 585 443
rect 367 417 585 425
rect 367 409 417 417
rect 367 375 375 409
rect 409 375 417 409
rect 535 409 585 417
rect 199 325 207 341
rect 73 307 207 325
rect 241 325 249 341
rect 367 341 417 375
rect 367 325 375 341
rect 241 307 375 325
rect 409 307 417 341
rect 30 291 417 307
rect 451 341 501 383
rect 535 375 543 409
rect 577 375 585 409
rect 535 359 585 375
rect 619 477 1005 493
rect 619 443 627 477
rect 661 459 795 477
rect 661 443 669 459
rect 619 409 669 443
rect 787 443 795 459
rect 829 459 963 477
rect 829 443 837 459
rect 787 427 837 443
rect 955 443 963 459
rect 997 443 1005 477
rect 955 427 1005 443
rect 1039 477 1089 493
rect 1039 459 1047 477
rect 1039 425 1041 459
rect 1081 443 1089 477
rect 1075 425 1089 443
rect 619 375 627 409
rect 661 375 669 409
rect 451 307 459 341
rect 493 325 501 341
rect 619 341 669 375
rect 703 409 753 425
rect 703 375 711 409
rect 745 393 753 409
rect 871 409 921 425
rect 871 393 879 409
rect 745 375 879 393
rect 913 391 921 409
rect 1123 391 1179 493
rect 913 375 1179 391
rect 703 357 1179 375
rect 619 325 627 341
rect 493 307 627 325
rect 661 307 669 341
rect 451 291 669 307
rect 703 289 1033 323
rect 703 257 737 289
rect 18 249 365 257
rect 18 215 99 249
rect 133 215 167 249
rect 201 215 235 249
rect 269 215 303 249
rect 337 215 365 249
rect 419 249 737 257
rect 999 257 1033 289
rect 419 215 435 249
rect 469 215 503 249
rect 537 215 737 249
rect 771 249 953 255
rect 771 215 823 249
rect 857 215 891 249
rect 925 215 953 249
rect 999 249 1083 257
rect 999 215 1015 249
rect 1049 215 1083 249
rect 1121 181 1179 357
rect 18 163 73 181
rect 18 129 39 163
rect 18 95 73 129
rect 18 61 39 95
rect 18 17 73 61
rect 107 163 1179 181
rect 107 129 123 163
rect 157 145 291 163
rect 157 129 173 145
rect 107 95 173 129
rect 275 129 291 145
rect 325 145 459 163
rect 325 129 341 145
rect 107 61 123 95
rect 157 61 173 95
rect 107 51 173 61
rect 207 95 241 111
rect 207 17 241 61
rect 275 95 341 129
rect 443 129 459 145
rect 493 145 627 163
rect 493 129 509 145
rect 275 61 291 95
rect 325 61 341 95
rect 275 51 341 61
rect 375 95 409 111
rect 375 17 409 61
rect 443 95 509 129
rect 611 129 627 145
rect 661 145 795 163
rect 661 129 677 145
rect 443 61 459 95
rect 493 61 509 95
rect 443 51 509 61
rect 543 95 577 111
rect 543 17 577 61
rect 611 95 677 129
rect 779 129 795 145
rect 829 145 963 163
rect 829 129 845 145
rect 611 61 627 95
rect 661 61 677 95
rect 611 51 677 61
rect 711 95 745 111
rect 711 17 745 61
rect 779 95 845 129
rect 947 129 963 145
rect 997 145 1179 163
rect 997 129 1013 145
rect 779 61 795 95
rect 829 61 845 95
rect 779 51 845 61
rect 879 95 913 111
rect 879 17 913 61
rect 947 95 1013 129
rect 947 61 963 95
rect 997 61 1013 95
rect 947 51 1013 61
rect 1047 95 1081 111
rect 1047 17 1081 61
rect 1121 51 1179 145
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 489 425 523 459
rect 1041 443 1047 459
rect 1047 443 1075 459
rect 1041 425 1075 443
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 477 459 536 467
rect 477 425 489 459
rect 523 456 536 459
rect 1029 459 1088 467
rect 1029 456 1041 459
rect 523 428 1041 456
rect 523 425 536 428
rect 477 413 536 425
rect 1029 425 1041 428
rect 1075 425 1088 459
rect 1029 413 1088 425
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 122 221 156 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 858 221 892 255 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 1133 289 1167 323 0 FreeSans 400 0 0 0 Y
port 8 nsew signal output
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nor3_4
rlabel metal1 s 0 -48 1196 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1196 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_END 2020068
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2010752
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 29.900 0.000 
<< end >>
