magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 1 21 1423 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 267 47 297 177
rect 351 47 381 177
rect 435 47 465 177
rect 519 47 549 177
rect 603 47 633 177
rect 687 47 717 177
rect 771 47 801 177
rect 855 47 885 177
rect 1043 47 1073 177
rect 1127 47 1157 177
rect 1211 47 1241 177
rect 1295 47 1325 177
<< scpmoshvt >>
rect 79 297 109 497
rect 267 297 297 497
rect 351 297 381 497
rect 435 297 465 497
rect 519 297 549 497
rect 603 297 633 497
rect 687 297 717 497
rect 771 297 801 497
rect 855 297 885 497
rect 1043 297 1073 497
rect 1127 297 1157 497
rect 1211 297 1241 497
rect 1295 297 1325 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 93 161 177
rect 109 59 119 93
rect 153 59 161 93
rect 109 47 161 59
rect 215 93 267 177
rect 215 59 223 93
rect 257 59 267 93
rect 215 47 267 59
rect 297 161 351 177
rect 297 127 307 161
rect 341 127 351 161
rect 297 47 351 127
rect 381 93 435 177
rect 381 59 391 93
rect 425 59 435 93
rect 381 47 435 59
rect 465 161 519 177
rect 465 127 475 161
rect 509 127 519 161
rect 465 47 519 127
rect 549 93 603 177
rect 549 59 559 93
rect 593 59 603 93
rect 549 47 603 59
rect 633 161 687 177
rect 633 127 643 161
rect 677 127 687 161
rect 633 47 687 127
rect 717 93 771 177
rect 717 59 727 93
rect 761 59 771 93
rect 717 47 771 59
rect 801 161 855 177
rect 801 127 811 161
rect 845 127 855 161
rect 801 47 855 127
rect 885 93 937 177
rect 885 59 895 93
rect 929 59 937 93
rect 885 47 937 59
rect 991 93 1043 177
rect 991 59 999 93
rect 1033 59 1043 93
rect 991 47 1043 59
rect 1073 161 1127 177
rect 1073 127 1083 161
rect 1117 127 1127 161
rect 1073 93 1127 127
rect 1073 59 1083 93
rect 1117 59 1127 93
rect 1073 47 1127 59
rect 1157 93 1211 177
rect 1157 59 1167 93
rect 1201 59 1211 93
rect 1157 47 1211 59
rect 1241 161 1295 177
rect 1241 127 1251 161
rect 1285 127 1295 161
rect 1241 93 1295 127
rect 1241 59 1251 93
rect 1285 59 1295 93
rect 1241 47 1295 59
rect 1325 161 1397 177
rect 1325 127 1351 161
rect 1385 127 1397 161
rect 1325 93 1397 127
rect 1325 59 1351 93
rect 1385 59 1397 93
rect 1325 47 1397 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 485 161 497
rect 109 451 119 485
rect 153 451 161 485
rect 109 417 161 451
rect 109 383 119 417
rect 153 383 161 417
rect 109 349 161 383
rect 109 315 119 349
rect 153 315 161 349
rect 109 297 161 315
rect 215 485 267 497
rect 215 451 223 485
rect 257 451 267 485
rect 215 417 267 451
rect 215 383 223 417
rect 257 383 267 417
rect 215 349 267 383
rect 215 315 223 349
rect 257 315 267 349
rect 215 297 267 315
rect 297 485 351 497
rect 297 451 307 485
rect 341 451 351 485
rect 297 417 351 451
rect 297 383 307 417
rect 341 383 351 417
rect 297 349 351 383
rect 297 315 307 349
rect 341 315 351 349
rect 297 297 351 315
rect 381 485 435 497
rect 381 451 391 485
rect 425 451 435 485
rect 381 417 435 451
rect 381 383 391 417
rect 425 383 435 417
rect 381 297 435 383
rect 465 485 519 497
rect 465 451 475 485
rect 509 451 519 485
rect 465 417 519 451
rect 465 383 475 417
rect 509 383 519 417
rect 465 349 519 383
rect 465 315 475 349
rect 509 315 519 349
rect 465 297 519 315
rect 549 485 603 497
rect 549 451 559 485
rect 593 451 603 485
rect 549 297 603 451
rect 633 485 687 497
rect 633 451 643 485
rect 677 451 687 485
rect 633 417 687 451
rect 633 383 643 417
rect 677 383 687 417
rect 633 349 687 383
rect 633 315 643 349
rect 677 315 687 349
rect 633 297 687 315
rect 717 485 771 497
rect 717 451 727 485
rect 761 451 771 485
rect 717 417 771 451
rect 717 383 727 417
rect 761 383 771 417
rect 717 297 771 383
rect 801 485 855 497
rect 801 451 811 485
rect 845 451 855 485
rect 801 417 855 451
rect 801 383 811 417
rect 845 383 855 417
rect 801 349 855 383
rect 801 315 811 349
rect 845 315 855 349
rect 801 297 855 315
rect 885 485 937 497
rect 885 451 895 485
rect 929 451 937 485
rect 885 417 937 451
rect 885 383 895 417
rect 929 383 937 417
rect 885 297 937 383
rect 991 485 1043 497
rect 991 451 999 485
rect 1033 451 1043 485
rect 991 417 1043 451
rect 991 383 999 417
rect 1033 383 1043 417
rect 991 297 1043 383
rect 1073 485 1127 497
rect 1073 451 1083 485
rect 1117 451 1127 485
rect 1073 417 1127 451
rect 1073 383 1083 417
rect 1117 383 1127 417
rect 1073 349 1127 383
rect 1073 315 1083 349
rect 1117 315 1127 349
rect 1073 297 1127 315
rect 1157 485 1211 497
rect 1157 451 1167 485
rect 1201 451 1211 485
rect 1157 417 1211 451
rect 1157 383 1167 417
rect 1201 383 1211 417
rect 1157 297 1211 383
rect 1241 485 1295 497
rect 1241 451 1251 485
rect 1285 451 1295 485
rect 1241 417 1295 451
rect 1241 383 1251 417
rect 1285 383 1295 417
rect 1241 349 1295 383
rect 1241 315 1251 349
rect 1285 315 1295 349
rect 1241 297 1295 315
rect 1325 485 1397 497
rect 1325 451 1351 485
rect 1385 451 1397 485
rect 1325 417 1397 451
rect 1325 383 1351 417
rect 1385 383 1397 417
rect 1325 349 1397 383
rect 1325 315 1351 349
rect 1385 315 1397 349
rect 1325 297 1397 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 119 59 153 93
rect 223 59 257 93
rect 307 127 341 161
rect 391 59 425 93
rect 475 127 509 161
rect 559 59 593 93
rect 643 127 677 161
rect 727 59 761 93
rect 811 127 845 161
rect 895 59 929 93
rect 999 59 1033 93
rect 1083 127 1117 161
rect 1083 59 1117 93
rect 1167 59 1201 93
rect 1251 127 1285 161
rect 1251 59 1285 93
rect 1351 127 1385 161
rect 1351 59 1385 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 451 153 485
rect 119 383 153 417
rect 119 315 153 349
rect 223 451 257 485
rect 223 383 257 417
rect 223 315 257 349
rect 307 451 341 485
rect 307 383 341 417
rect 307 315 341 349
rect 391 451 425 485
rect 391 383 425 417
rect 475 451 509 485
rect 475 383 509 417
rect 475 315 509 349
rect 559 451 593 485
rect 643 451 677 485
rect 643 383 677 417
rect 643 315 677 349
rect 727 451 761 485
rect 727 383 761 417
rect 811 451 845 485
rect 811 383 845 417
rect 811 315 845 349
rect 895 451 929 485
rect 895 383 929 417
rect 999 451 1033 485
rect 999 383 1033 417
rect 1083 451 1117 485
rect 1083 383 1117 417
rect 1083 315 1117 349
rect 1167 451 1201 485
rect 1167 383 1201 417
rect 1251 451 1285 485
rect 1251 383 1285 417
rect 1251 315 1285 349
rect 1351 451 1385 485
rect 1351 383 1385 417
rect 1351 315 1385 349
<< poly >>
rect 79 497 109 523
rect 267 497 297 523
rect 351 497 381 523
rect 435 497 465 523
rect 519 497 549 523
rect 603 497 633 523
rect 687 497 717 523
rect 771 497 801 523
rect 855 497 885 523
rect 1043 497 1073 523
rect 1127 497 1157 523
rect 1211 497 1241 523
rect 1295 497 1325 523
rect 79 261 109 297
rect 79 249 152 261
rect 267 259 297 297
rect 351 259 381 297
rect 435 259 465 297
rect 519 259 549 297
rect 79 215 102 249
rect 136 215 152 249
rect 79 203 152 215
rect 201 249 549 259
rect 201 215 217 249
rect 251 215 307 249
rect 341 215 391 249
rect 425 215 475 249
rect 509 215 549 249
rect 201 205 549 215
rect 79 177 109 203
rect 267 177 297 205
rect 351 177 381 205
rect 435 177 465 205
rect 519 177 549 205
rect 603 259 633 297
rect 687 259 717 297
rect 771 259 801 297
rect 855 259 885 297
rect 1043 259 1073 297
rect 1127 259 1157 297
rect 1211 259 1241 297
rect 1295 259 1325 297
rect 603 249 885 259
rect 603 215 670 249
rect 704 215 806 249
rect 840 215 885 249
rect 603 205 885 215
rect 977 249 1325 259
rect 977 215 993 249
rect 1027 215 1083 249
rect 1117 215 1167 249
rect 1201 215 1250 249
rect 1284 215 1325 249
rect 977 205 1325 215
rect 603 177 633 205
rect 687 177 717 205
rect 771 177 801 205
rect 855 177 885 205
rect 1043 177 1073 205
rect 1127 177 1157 205
rect 1211 177 1241 205
rect 1295 177 1325 205
rect 79 21 109 47
rect 267 21 297 47
rect 351 21 381 47
rect 435 21 465 47
rect 519 21 549 47
rect 603 21 633 47
rect 687 21 717 47
rect 771 21 801 47
rect 855 21 885 47
rect 1043 21 1073 47
rect 1127 21 1157 47
rect 1211 21 1241 47
rect 1295 21 1325 47
<< polycont >>
rect 102 215 136 249
rect 217 215 251 249
rect 307 215 341 249
rect 391 215 425 249
rect 475 215 509 249
rect 670 215 704 249
rect 806 215 840 249
rect 993 215 1027 249
rect 1083 215 1117 249
rect 1167 215 1201 249
rect 1250 215 1284 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 17 485 85 493
rect 17 451 35 485
rect 69 451 85 485
rect 17 417 85 451
rect 17 383 35 417
rect 69 383 85 417
rect 17 349 85 383
rect 17 315 35 349
rect 69 315 85 349
rect 17 289 85 315
rect 119 485 257 527
rect 153 451 223 485
rect 119 417 257 451
rect 153 383 223 417
rect 119 349 257 383
rect 153 315 223 349
rect 119 289 257 315
rect 291 485 357 493
rect 291 451 307 485
rect 341 451 357 485
rect 291 417 357 451
rect 291 383 307 417
rect 341 383 357 417
rect 291 349 357 383
rect 391 485 425 527
rect 391 417 425 451
rect 391 367 425 383
rect 459 485 525 493
rect 459 451 475 485
rect 509 451 525 485
rect 459 417 525 451
rect 559 485 593 527
rect 559 435 593 451
rect 627 485 693 493
rect 627 451 643 485
rect 677 451 693 485
rect 459 383 475 417
rect 509 401 525 417
rect 627 417 693 451
rect 627 401 643 417
rect 509 383 643 401
rect 677 383 693 417
rect 291 315 307 349
rect 341 333 357 349
rect 459 349 693 383
rect 727 485 761 527
rect 727 417 761 451
rect 727 367 761 383
rect 795 485 861 493
rect 795 451 811 485
rect 845 451 861 485
rect 795 417 861 451
rect 795 383 811 417
rect 845 383 861 417
rect 459 333 475 349
rect 341 315 475 333
rect 509 315 643 349
rect 677 333 693 349
rect 795 349 861 383
rect 895 485 1033 527
rect 929 451 999 485
rect 895 417 1033 451
rect 929 383 999 417
rect 895 367 1033 383
rect 1067 485 1133 493
rect 1067 451 1083 485
rect 1117 451 1133 485
rect 1067 417 1133 451
rect 1067 383 1083 417
rect 1117 383 1133 417
rect 795 333 811 349
rect 677 315 811 333
rect 845 333 861 349
rect 1067 349 1133 383
rect 1167 485 1201 527
rect 1167 417 1201 451
rect 1167 367 1201 383
rect 1235 485 1301 493
rect 1235 451 1251 485
rect 1285 451 1301 485
rect 1235 417 1301 451
rect 1235 383 1251 417
rect 1285 383 1301 417
rect 1067 333 1083 349
rect 845 315 1083 333
rect 1117 333 1133 349
rect 1235 349 1301 383
rect 1235 333 1251 349
rect 1117 315 1251 333
rect 1285 315 1301 349
rect 291 289 1301 315
rect 1335 485 1401 527
rect 1335 451 1351 485
rect 1385 451 1401 485
rect 1335 417 1401 451
rect 1335 383 1351 417
rect 1385 383 1401 417
rect 1335 349 1401 383
rect 1335 315 1351 349
rect 1385 315 1401 349
rect 1335 289 1401 315
rect 17 181 52 289
rect 86 249 156 255
rect 86 215 102 249
rect 136 215 156 249
rect 201 249 525 255
rect 201 215 217 249
rect 251 215 307 249
rect 341 215 391 249
rect 425 215 475 249
rect 509 215 525 249
rect 559 215 620 289
rect 654 249 896 255
rect 654 215 670 249
rect 704 215 806 249
rect 840 215 896 249
rect 958 249 1300 255
rect 958 215 993 249
rect 1027 215 1083 249
rect 1117 215 1167 249
rect 1201 215 1250 249
rect 1284 215 1300 249
rect 201 181 257 215
rect 559 181 593 215
rect 17 161 257 181
rect 17 127 35 161
rect 69 143 257 161
rect 291 161 593 181
rect 69 127 85 143
rect 291 127 307 161
rect 341 127 475 161
rect 509 127 593 161
rect 627 161 1301 181
rect 627 127 643 161
rect 677 127 811 161
rect 845 143 1083 161
rect 845 127 945 143
rect 1067 127 1083 143
rect 1117 143 1251 161
rect 1117 127 1133 143
rect 17 93 85 127
rect 17 59 35 93
rect 69 59 85 93
rect 17 51 85 59
rect 119 93 169 109
rect 983 93 1033 109
rect 153 59 169 93
rect 119 17 169 59
rect 207 59 223 93
rect 257 59 391 93
rect 425 59 559 93
rect 593 59 727 93
rect 761 59 895 93
rect 929 59 945 93
rect 207 51 945 59
rect 983 59 999 93
rect 983 17 1033 59
rect 1067 93 1133 127
rect 1235 127 1251 143
rect 1285 127 1301 161
rect 1067 59 1083 93
rect 1117 59 1133 93
rect 1067 51 1133 59
rect 1167 93 1201 109
rect 1167 17 1201 59
rect 1235 93 1301 127
rect 1235 59 1251 93
rect 1285 59 1301 93
rect 1235 51 1301 59
rect 1335 161 1401 181
rect 1335 127 1351 161
rect 1385 127 1401 161
rect 1335 93 1401 127
rect 1335 59 1351 93
rect 1385 59 1401 93
rect 1335 17 1401 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 586 221 620 255 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 586 357 620 391 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 862 221 896 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 770 221 804 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 678 221 712 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 958 221 992 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 1050 221 1084 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 1142 221 1176 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 1234 221 1268 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 586 289 620 323 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nand3b_4
rlabel metal1 s 0 -48 1472 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1472 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1472 544
string GDS_END 1867596
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1855810
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 36.800 0.000 
<< end >>
