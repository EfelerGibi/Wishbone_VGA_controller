magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< poly >>
rect 297 435 327 648
rect 921 559 951 648
rect 903 543 969 559
rect 903 509 919 543
rect 953 509 969 543
rect 903 493 969 509
rect 1545 435 1575 648
rect 2169 559 2199 648
rect 2151 543 2217 559
rect 2151 509 2167 543
rect 2201 509 2217 543
rect 2151 493 2217 509
rect 2793 435 2823 648
rect 3417 559 3447 648
rect 3399 543 3465 559
rect 3399 509 3415 543
rect 3449 509 3465 543
rect 3399 493 3465 509
rect 4041 435 4071 648
rect 4665 559 4695 648
rect 4647 543 4713 559
rect 4647 509 4663 543
rect 4697 509 4713 543
rect 4647 493 4713 509
rect 5289 435 5319 648
rect 5913 559 5943 648
rect 5895 543 5961 559
rect 5895 509 5911 543
rect 5945 509 5961 543
rect 5895 493 5961 509
rect 6537 435 6567 648
rect 7161 559 7191 648
rect 7143 543 7209 559
rect 7143 509 7159 543
rect 7193 509 7209 543
rect 7143 493 7209 509
rect 7785 435 7815 648
rect 8409 559 8439 648
rect 8391 543 8457 559
rect 8391 509 8407 543
rect 8441 509 8457 543
rect 8391 493 8457 509
rect 9033 435 9063 648
rect 9657 559 9687 648
rect 9639 543 9705 559
rect 9639 509 9655 543
rect 9689 509 9705 543
rect 9639 493 9705 509
rect 10281 435 10311 648
rect 10905 559 10935 648
rect 10887 543 10953 559
rect 10887 509 10903 543
rect 10937 509 10953 543
rect 10887 493 10953 509
rect 11529 435 11559 648
rect 12153 559 12183 648
rect 12135 543 12201 559
rect 12135 509 12151 543
rect 12185 509 12201 543
rect 12135 493 12201 509
rect 12777 435 12807 648
rect 13401 559 13431 648
rect 13383 543 13449 559
rect 13383 509 13399 543
rect 13433 509 13449 543
rect 13383 493 13449 509
rect 14025 435 14055 648
rect 14649 559 14679 648
rect 14631 543 14697 559
rect 14631 509 14647 543
rect 14681 509 14697 543
rect 14631 493 14697 509
rect 15273 435 15303 648
rect 15897 559 15927 648
rect 15879 543 15945 559
rect 15879 509 15895 543
rect 15929 509 15945 543
rect 15879 493 15945 509
rect 16521 435 16551 648
rect 17145 559 17175 648
rect 17127 543 17193 559
rect 17127 509 17143 543
rect 17177 509 17193 543
rect 17127 493 17193 509
rect 17769 435 17799 648
rect 18393 559 18423 648
rect 18375 543 18441 559
rect 18375 509 18391 543
rect 18425 509 18441 543
rect 18375 493 18441 509
rect 19017 435 19047 648
rect 19641 559 19671 648
rect 19623 543 19689 559
rect 19623 509 19639 543
rect 19673 509 19689 543
rect 19623 493 19689 509
rect 20265 435 20295 648
rect 20889 559 20919 648
rect 20871 543 20937 559
rect 20871 509 20887 543
rect 20921 509 20937 543
rect 20871 493 20937 509
rect 21513 435 21543 648
rect 22137 559 22167 648
rect 22119 543 22185 559
rect 22119 509 22135 543
rect 22169 509 22185 543
rect 22119 493 22185 509
rect 22761 435 22791 648
rect 23385 559 23415 648
rect 23367 543 23433 559
rect 23367 509 23383 543
rect 23417 509 23433 543
rect 23367 493 23433 509
rect 24009 435 24039 648
rect 24633 559 24663 648
rect 24615 543 24681 559
rect 24615 509 24631 543
rect 24665 509 24681 543
rect 24615 493 24681 509
rect 25257 435 25287 648
rect 25881 559 25911 648
rect 25863 543 25929 559
rect 25863 509 25879 543
rect 25913 509 25929 543
rect 25863 493 25929 509
rect 26505 435 26535 648
rect 27129 559 27159 648
rect 27111 543 27177 559
rect 27111 509 27127 543
rect 27161 509 27177 543
rect 27111 493 27177 509
rect 27753 435 27783 648
rect 28377 559 28407 648
rect 28359 543 28425 559
rect 28359 509 28375 543
rect 28409 509 28425 543
rect 28359 493 28425 509
rect 29001 435 29031 648
rect 29625 559 29655 648
rect 29607 543 29673 559
rect 29607 509 29623 543
rect 29657 509 29673 543
rect 29607 493 29673 509
rect 30249 435 30279 648
rect 30873 559 30903 648
rect 30855 543 30921 559
rect 30855 509 30871 543
rect 30905 509 30921 543
rect 30855 493 30921 509
rect 31497 435 31527 648
rect 32121 559 32151 648
rect 32103 543 32169 559
rect 32103 509 32119 543
rect 32153 509 32169 543
rect 32103 493 32169 509
rect 32745 435 32775 648
rect 33369 559 33399 648
rect 33351 543 33417 559
rect 33351 509 33367 543
rect 33401 509 33417 543
rect 33351 493 33417 509
rect 33993 435 34023 648
rect 34617 559 34647 648
rect 34599 543 34665 559
rect 34599 509 34615 543
rect 34649 509 34665 543
rect 34599 493 34665 509
rect 35241 435 35271 648
rect 35865 559 35895 648
rect 35847 543 35913 559
rect 35847 509 35863 543
rect 35897 509 35913 543
rect 35847 493 35913 509
rect 36489 435 36519 648
rect 37113 559 37143 648
rect 37095 543 37161 559
rect 37095 509 37111 543
rect 37145 509 37161 543
rect 37095 493 37161 509
rect 37737 435 37767 648
rect 38361 559 38391 648
rect 38343 543 38409 559
rect 38343 509 38359 543
rect 38393 509 38409 543
rect 38343 493 38409 509
rect 38985 435 39015 648
rect 39609 559 39639 648
rect 39591 543 39657 559
rect 39591 509 39607 543
rect 39641 509 39657 543
rect 39591 493 39657 509
rect 279 419 345 435
rect 279 385 295 419
rect 329 385 345 419
rect 279 369 345 385
rect 1527 419 1593 435
rect 1527 385 1543 419
rect 1577 385 1593 419
rect 1527 369 1593 385
rect 2775 419 2841 435
rect 2775 385 2791 419
rect 2825 385 2841 419
rect 2775 369 2841 385
rect 4023 419 4089 435
rect 4023 385 4039 419
rect 4073 385 4089 419
rect 4023 369 4089 385
rect 5271 419 5337 435
rect 5271 385 5287 419
rect 5321 385 5337 419
rect 5271 369 5337 385
rect 6519 419 6585 435
rect 6519 385 6535 419
rect 6569 385 6585 419
rect 6519 369 6585 385
rect 7767 419 7833 435
rect 7767 385 7783 419
rect 7817 385 7833 419
rect 7767 369 7833 385
rect 9015 419 9081 435
rect 9015 385 9031 419
rect 9065 385 9081 419
rect 9015 369 9081 385
rect 10263 419 10329 435
rect 10263 385 10279 419
rect 10313 385 10329 419
rect 10263 369 10329 385
rect 11511 419 11577 435
rect 11511 385 11527 419
rect 11561 385 11577 419
rect 11511 369 11577 385
rect 12759 419 12825 435
rect 12759 385 12775 419
rect 12809 385 12825 419
rect 12759 369 12825 385
rect 14007 419 14073 435
rect 14007 385 14023 419
rect 14057 385 14073 419
rect 14007 369 14073 385
rect 15255 419 15321 435
rect 15255 385 15271 419
rect 15305 385 15321 419
rect 15255 369 15321 385
rect 16503 419 16569 435
rect 16503 385 16519 419
rect 16553 385 16569 419
rect 16503 369 16569 385
rect 17751 419 17817 435
rect 17751 385 17767 419
rect 17801 385 17817 419
rect 17751 369 17817 385
rect 18999 419 19065 435
rect 18999 385 19015 419
rect 19049 385 19065 419
rect 18999 369 19065 385
rect 20247 419 20313 435
rect 20247 385 20263 419
rect 20297 385 20313 419
rect 20247 369 20313 385
rect 21495 419 21561 435
rect 21495 385 21511 419
rect 21545 385 21561 419
rect 21495 369 21561 385
rect 22743 419 22809 435
rect 22743 385 22759 419
rect 22793 385 22809 419
rect 22743 369 22809 385
rect 23991 419 24057 435
rect 23991 385 24007 419
rect 24041 385 24057 419
rect 23991 369 24057 385
rect 25239 419 25305 435
rect 25239 385 25255 419
rect 25289 385 25305 419
rect 25239 369 25305 385
rect 26487 419 26553 435
rect 26487 385 26503 419
rect 26537 385 26553 419
rect 26487 369 26553 385
rect 27735 419 27801 435
rect 27735 385 27751 419
rect 27785 385 27801 419
rect 27735 369 27801 385
rect 28983 419 29049 435
rect 28983 385 28999 419
rect 29033 385 29049 419
rect 28983 369 29049 385
rect 30231 419 30297 435
rect 30231 385 30247 419
rect 30281 385 30297 419
rect 30231 369 30297 385
rect 31479 419 31545 435
rect 31479 385 31495 419
rect 31529 385 31545 419
rect 31479 369 31545 385
rect 32727 419 32793 435
rect 32727 385 32743 419
rect 32777 385 32793 419
rect 32727 369 32793 385
rect 33975 419 34041 435
rect 33975 385 33991 419
rect 34025 385 34041 419
rect 33975 369 34041 385
rect 35223 419 35289 435
rect 35223 385 35239 419
rect 35273 385 35289 419
rect 35223 369 35289 385
rect 36471 419 36537 435
rect 36471 385 36487 419
rect 36521 385 36537 419
rect 36471 369 36537 385
rect 37719 419 37785 435
rect 37719 385 37735 419
rect 37769 385 37785 419
rect 37719 369 37785 385
rect 38967 419 39033 435
rect 38967 385 38983 419
rect 39017 385 39033 419
rect 38967 369 39033 385
<< polycont >>
rect 919 509 953 543
rect 2167 509 2201 543
rect 3415 509 3449 543
rect 4663 509 4697 543
rect 5911 509 5945 543
rect 7159 509 7193 543
rect 8407 509 8441 543
rect 9655 509 9689 543
rect 10903 509 10937 543
rect 12151 509 12185 543
rect 13399 509 13433 543
rect 14647 509 14681 543
rect 15895 509 15929 543
rect 17143 509 17177 543
rect 18391 509 18425 543
rect 19639 509 19673 543
rect 20887 509 20921 543
rect 22135 509 22169 543
rect 23383 509 23417 543
rect 24631 509 24665 543
rect 25879 509 25913 543
rect 27127 509 27161 543
rect 28375 509 28409 543
rect 29623 509 29657 543
rect 30871 509 30905 543
rect 32119 509 32153 543
rect 33367 509 33401 543
rect 34615 509 34649 543
rect 35863 509 35897 543
rect 37111 509 37145 543
rect 38359 509 38393 543
rect 39607 509 39641 543
rect 295 385 329 419
rect 1543 385 1577 419
rect 2791 385 2825 419
rect 4039 385 4073 419
rect 5287 385 5321 419
rect 6535 385 6569 419
rect 7783 385 7817 419
rect 9031 385 9065 419
rect 10279 385 10313 419
rect 11527 385 11561 419
rect 12775 385 12809 419
rect 14023 385 14057 419
rect 15271 385 15305 419
rect 16519 385 16553 419
rect 17767 385 17801 419
rect 19015 385 19049 419
rect 20263 385 20297 419
rect 21511 385 21545 419
rect 22759 385 22793 419
rect 24007 385 24041 419
rect 25255 385 25289 419
rect 26503 385 26537 419
rect 27751 385 27785 419
rect 28999 385 29033 419
rect 30247 385 30281 419
rect 31495 385 31529 419
rect 32743 385 32777 419
rect 33991 385 34025 419
rect 35239 385 35273 419
rect 36487 385 36521 419
rect 37735 385 37769 419
rect 38983 385 39017 419
<< locali >>
rect 919 543 953 559
rect 919 493 953 509
rect 2167 543 2201 559
rect 2167 493 2201 509
rect 3415 543 3449 559
rect 3415 493 3449 509
rect 4663 543 4697 559
rect 4663 493 4697 509
rect 5911 543 5945 559
rect 5911 493 5945 509
rect 7159 543 7193 559
rect 7159 493 7193 509
rect 8407 543 8441 559
rect 8407 493 8441 509
rect 9655 543 9689 559
rect 9655 493 9689 509
rect 10903 543 10937 559
rect 10903 493 10937 509
rect 12151 543 12185 559
rect 12151 493 12185 509
rect 13399 543 13433 559
rect 13399 493 13433 509
rect 14647 543 14681 559
rect 14647 493 14681 509
rect 15895 543 15929 559
rect 15895 493 15929 509
rect 17143 543 17177 559
rect 17143 493 17177 509
rect 18391 543 18425 559
rect 18391 493 18425 509
rect 19639 543 19673 559
rect 19639 493 19673 509
rect 20887 543 20921 559
rect 20887 493 20921 509
rect 22135 543 22169 559
rect 22135 493 22169 509
rect 23383 543 23417 559
rect 23383 493 23417 509
rect 24631 543 24665 559
rect 24631 493 24665 509
rect 25879 543 25913 559
rect 25879 493 25913 509
rect 27127 543 27161 559
rect 27127 493 27161 509
rect 28375 543 28409 559
rect 28375 493 28409 509
rect 29623 543 29657 559
rect 29623 493 29657 509
rect 30871 543 30905 559
rect 30871 493 30905 509
rect 32119 543 32153 559
rect 32119 493 32153 509
rect 33367 543 33401 559
rect 33367 493 33401 509
rect 34615 543 34649 559
rect 34615 493 34649 509
rect 35863 543 35897 559
rect 35863 493 35897 509
rect 37111 543 37145 559
rect 37111 493 37145 509
rect 38359 543 38393 559
rect 38359 493 38393 509
rect 39607 543 39641 559
rect 39607 493 39641 509
rect 295 419 329 435
rect 295 369 329 385
rect 1543 419 1577 435
rect 1543 369 1577 385
rect 2791 419 2825 435
rect 2791 369 2825 385
rect 4039 419 4073 435
rect 4039 369 4073 385
rect 5287 419 5321 435
rect 5287 369 5321 385
rect 6535 419 6569 435
rect 6535 369 6569 385
rect 7783 419 7817 435
rect 7783 369 7817 385
rect 9031 419 9065 435
rect 9031 369 9065 385
rect 10279 419 10313 435
rect 10279 369 10313 385
rect 11527 419 11561 435
rect 11527 369 11561 385
rect 12775 419 12809 435
rect 12775 369 12809 385
rect 14023 419 14057 435
rect 14023 369 14057 385
rect 15271 419 15305 435
rect 15271 369 15305 385
rect 16519 419 16553 435
rect 16519 369 16553 385
rect 17767 419 17801 435
rect 17767 369 17801 385
rect 19015 419 19049 435
rect 19015 369 19049 385
rect 20263 419 20297 435
rect 20263 369 20297 385
rect 21511 419 21545 435
rect 21511 369 21545 385
rect 22759 419 22793 435
rect 22759 369 22793 385
rect 24007 419 24041 435
rect 24007 369 24041 385
rect 25255 419 25289 435
rect 25255 369 25289 385
rect 26503 419 26537 435
rect 26503 369 26537 385
rect 27751 419 27785 435
rect 27751 369 27785 385
rect 28999 419 29033 435
rect 28999 369 29033 385
rect 30247 419 30281 435
rect 30247 369 30281 385
rect 31495 419 31529 435
rect 31495 369 31529 385
rect 32743 419 32777 435
rect 32743 369 32777 385
rect 33991 419 34025 435
rect 33991 369 34025 385
rect 35239 419 35273 435
rect 35239 369 35273 385
rect 36487 419 36521 435
rect 36487 369 36521 385
rect 37735 419 37769 435
rect 37735 369 37769 385
rect 38983 419 39017 435
rect 38983 369 39017 385
<< viali >>
rect 919 509 953 543
rect 2167 509 2201 543
rect 3415 509 3449 543
rect 4663 509 4697 543
rect 5911 509 5945 543
rect 7159 509 7193 543
rect 8407 509 8441 543
rect 9655 509 9689 543
rect 10903 509 10937 543
rect 12151 509 12185 543
rect 13399 509 13433 543
rect 14647 509 14681 543
rect 15895 509 15929 543
rect 17143 509 17177 543
rect 18391 509 18425 543
rect 19639 509 19673 543
rect 20887 509 20921 543
rect 22135 509 22169 543
rect 23383 509 23417 543
rect 24631 509 24665 543
rect 25879 509 25913 543
rect 27127 509 27161 543
rect 28375 509 28409 543
rect 29623 509 29657 543
rect 30871 509 30905 543
rect 32119 509 32153 543
rect 33367 509 33401 543
rect 34615 509 34649 543
rect 35863 509 35897 543
rect 37111 509 37145 543
rect 38359 509 38393 543
rect 39607 509 39641 543
rect 295 385 329 419
rect 1543 385 1577 419
rect 2791 385 2825 419
rect 4039 385 4073 419
rect 5287 385 5321 419
rect 6535 385 6569 419
rect 7783 385 7817 419
rect 9031 385 9065 419
rect 10279 385 10313 419
rect 11527 385 11561 419
rect 12775 385 12809 419
rect 14023 385 14057 419
rect 15271 385 15305 419
rect 16519 385 16553 419
rect 17767 385 17801 419
rect 19015 385 19049 419
rect 20263 385 20297 419
rect 21511 385 21545 419
rect 22759 385 22793 419
rect 24007 385 24041 419
rect 25255 385 25289 419
rect 26503 385 26537 419
rect 27751 385 27785 419
rect 28999 385 29033 419
rect 30247 385 30281 419
rect 31495 385 31529 419
rect 32743 385 32777 419
rect 33991 385 34025 419
rect 35239 385 35273 419
rect 36487 385 36521 419
rect 37735 385 37769 419
rect 38983 385 39017 419
<< metal1 >>
rect 80 1928 108 1984
rect 544 1928 572 1984
rect 676 1928 704 1984
rect 1140 1928 1168 1984
rect 1328 1928 1356 1984
rect 1792 1928 1820 1984
rect 1924 1928 1952 1984
rect 2388 1928 2416 1984
rect 2576 1928 2604 1984
rect 3040 1928 3068 1984
rect 3172 1928 3200 1984
rect 3636 1928 3664 1984
rect 3824 1928 3852 1984
rect 4288 1928 4316 1984
rect 4420 1928 4448 1984
rect 4884 1928 4912 1984
rect 5072 1928 5100 1984
rect 5536 1928 5564 1984
rect 5668 1928 5696 1984
rect 6132 1928 6160 1984
rect 6320 1928 6348 1984
rect 6784 1928 6812 1984
rect 6916 1928 6944 1984
rect 7380 1928 7408 1984
rect 7568 1928 7596 1984
rect 8032 1928 8060 1984
rect 8164 1928 8192 1984
rect 8628 1928 8656 1984
rect 8816 1928 8844 1984
rect 9280 1928 9308 1984
rect 9412 1928 9440 1984
rect 9876 1928 9904 1984
rect 10064 1928 10092 1984
rect 10528 1928 10556 1984
rect 10660 1928 10688 1984
rect 11124 1928 11152 1984
rect 11312 1928 11340 1984
rect 11776 1928 11804 1984
rect 11908 1928 11936 1984
rect 12372 1928 12400 1984
rect 12560 1928 12588 1984
rect 13024 1928 13052 1984
rect 13156 1928 13184 1984
rect 13620 1928 13648 1984
rect 13808 1928 13836 1984
rect 14272 1928 14300 1984
rect 14404 1928 14432 1984
rect 14868 1928 14896 1984
rect 15056 1928 15084 1984
rect 15520 1928 15548 1984
rect 15652 1928 15680 1984
rect 16116 1928 16144 1984
rect 16304 1928 16332 1984
rect 16768 1928 16796 1984
rect 16900 1928 16928 1984
rect 17364 1928 17392 1984
rect 17552 1928 17580 1984
rect 18016 1928 18044 1984
rect 18148 1928 18176 1984
rect 18612 1928 18640 1984
rect 18800 1928 18828 1984
rect 19264 1928 19292 1984
rect 19396 1928 19424 1984
rect 19860 1928 19888 1984
rect 20048 1928 20076 1984
rect 20512 1928 20540 1984
rect 20644 1928 20672 1984
rect 21108 1928 21136 1984
rect 21296 1928 21324 1984
rect 21760 1928 21788 1984
rect 21892 1928 21920 1984
rect 22356 1928 22384 1984
rect 22544 1928 22572 1984
rect 23008 1928 23036 1984
rect 23140 1928 23168 1984
rect 23604 1928 23632 1984
rect 23792 1928 23820 1984
rect 24256 1928 24284 1984
rect 24388 1928 24416 1984
rect 24852 1928 24880 1984
rect 25040 1928 25068 1984
rect 25504 1928 25532 1984
rect 25636 1928 25664 1984
rect 26100 1928 26128 1984
rect 26288 1928 26316 1984
rect 26752 1928 26780 1984
rect 26884 1928 26912 1984
rect 27348 1928 27376 1984
rect 27536 1928 27564 1984
rect 28000 1928 28028 1984
rect 28132 1928 28160 1984
rect 28596 1928 28624 1984
rect 28784 1928 28812 1984
rect 29248 1928 29276 1984
rect 29380 1928 29408 1984
rect 29844 1928 29872 1984
rect 30032 1928 30060 1984
rect 30496 1928 30524 1984
rect 30628 1928 30656 1984
rect 31092 1928 31120 1984
rect 31280 1928 31308 1984
rect 31744 1928 31772 1984
rect 31876 1928 31904 1984
rect 32340 1928 32368 1984
rect 32528 1928 32556 1984
rect 32992 1928 33020 1984
rect 33124 1928 33152 1984
rect 33588 1928 33616 1984
rect 33776 1928 33804 1984
rect 34240 1928 34268 1984
rect 34372 1928 34400 1984
rect 34836 1928 34864 1984
rect 35024 1928 35052 1984
rect 35488 1928 35516 1984
rect 35620 1928 35648 1984
rect 36084 1928 36112 1984
rect 36272 1928 36300 1984
rect 36736 1928 36764 1984
rect 36868 1928 36896 1984
rect 37332 1928 37360 1984
rect 37520 1928 37548 1984
rect 37984 1928 38012 1984
rect 38116 1928 38144 1984
rect 38580 1928 38608 1984
rect 38768 1928 38796 1984
rect 39232 1928 39260 1984
rect 39364 1928 39392 1984
rect 39828 1928 39856 1984
rect 80 274 108 620
rect 280 376 286 428
rect 338 376 344 428
rect 62 222 68 274
rect 120 222 126 274
rect 544 150 572 620
rect 676 150 704 620
rect 904 500 910 552
rect 962 500 968 552
rect 1140 274 1168 620
rect 1328 274 1356 620
rect 1528 376 1534 428
rect 1586 376 1592 428
rect 1122 222 1128 274
rect 1180 222 1186 274
rect 1310 222 1316 274
rect 1368 222 1374 274
rect 1792 150 1820 620
rect 1924 150 1952 620
rect 2152 500 2158 552
rect 2210 500 2216 552
rect 2388 274 2416 620
rect 2576 274 2604 620
rect 2776 376 2782 428
rect 2834 376 2840 428
rect 2370 222 2376 274
rect 2428 222 2434 274
rect 2558 222 2564 274
rect 2616 222 2622 274
rect 3040 150 3068 620
rect 3172 150 3200 620
rect 3400 500 3406 552
rect 3458 500 3464 552
rect 3636 274 3664 620
rect 3824 274 3852 620
rect 4024 376 4030 428
rect 4082 376 4088 428
rect 3618 222 3624 274
rect 3676 222 3682 274
rect 3806 222 3812 274
rect 3864 222 3870 274
rect 4288 150 4316 620
rect 4420 150 4448 620
rect 4648 500 4654 552
rect 4706 500 4712 552
rect 4884 274 4912 620
rect 5072 274 5100 620
rect 5272 376 5278 428
rect 5330 376 5336 428
rect 4866 222 4872 274
rect 4924 222 4930 274
rect 5054 222 5060 274
rect 5112 222 5118 274
rect 5536 150 5564 620
rect 5668 150 5696 620
rect 5896 500 5902 552
rect 5954 500 5960 552
rect 6132 274 6160 620
rect 6320 274 6348 620
rect 6520 376 6526 428
rect 6578 376 6584 428
rect 6114 222 6120 274
rect 6172 222 6178 274
rect 6302 222 6308 274
rect 6360 222 6366 274
rect 6784 150 6812 620
rect 6916 150 6944 620
rect 7144 500 7150 552
rect 7202 500 7208 552
rect 7380 274 7408 620
rect 7568 274 7596 620
rect 7768 376 7774 428
rect 7826 376 7832 428
rect 7362 222 7368 274
rect 7420 222 7426 274
rect 7550 222 7556 274
rect 7608 222 7614 274
rect 8032 150 8060 620
rect 8164 150 8192 620
rect 8392 500 8398 552
rect 8450 500 8456 552
rect 8628 274 8656 620
rect 8816 274 8844 620
rect 9016 376 9022 428
rect 9074 376 9080 428
rect 8610 222 8616 274
rect 8668 222 8674 274
rect 8798 222 8804 274
rect 8856 222 8862 274
rect 9280 150 9308 620
rect 9412 150 9440 620
rect 9640 500 9646 552
rect 9698 500 9704 552
rect 9876 274 9904 620
rect 10064 274 10092 620
rect 10264 376 10270 428
rect 10322 376 10328 428
rect 9858 222 9864 274
rect 9916 222 9922 274
rect 10046 222 10052 274
rect 10104 222 10110 274
rect 10528 150 10556 620
rect 10660 150 10688 620
rect 10888 500 10894 552
rect 10946 500 10952 552
rect 11124 274 11152 620
rect 11312 274 11340 620
rect 11512 376 11518 428
rect 11570 376 11576 428
rect 11106 222 11112 274
rect 11164 222 11170 274
rect 11294 222 11300 274
rect 11352 222 11358 274
rect 11776 150 11804 620
rect 11908 150 11936 620
rect 12136 500 12142 552
rect 12194 500 12200 552
rect 12372 274 12400 620
rect 12560 274 12588 620
rect 12760 376 12766 428
rect 12818 376 12824 428
rect 12354 222 12360 274
rect 12412 222 12418 274
rect 12542 222 12548 274
rect 12600 222 12606 274
rect 13024 150 13052 620
rect 13156 150 13184 620
rect 13384 500 13390 552
rect 13442 500 13448 552
rect 13620 274 13648 620
rect 13808 274 13836 620
rect 14008 376 14014 428
rect 14066 376 14072 428
rect 13602 222 13608 274
rect 13660 222 13666 274
rect 13790 222 13796 274
rect 13848 222 13854 274
rect 14272 150 14300 620
rect 14404 150 14432 620
rect 14632 500 14638 552
rect 14690 500 14696 552
rect 14868 274 14896 620
rect 15056 274 15084 620
rect 15256 376 15262 428
rect 15314 376 15320 428
rect 14850 222 14856 274
rect 14908 222 14914 274
rect 15038 222 15044 274
rect 15096 222 15102 274
rect 15520 150 15548 620
rect 15652 150 15680 620
rect 15880 500 15886 552
rect 15938 500 15944 552
rect 16116 274 16144 620
rect 16304 274 16332 620
rect 16504 376 16510 428
rect 16562 376 16568 428
rect 16098 222 16104 274
rect 16156 222 16162 274
rect 16286 222 16292 274
rect 16344 222 16350 274
rect 16768 150 16796 620
rect 16900 150 16928 620
rect 17128 500 17134 552
rect 17186 500 17192 552
rect 17364 274 17392 620
rect 17552 274 17580 620
rect 17752 376 17758 428
rect 17810 376 17816 428
rect 17346 222 17352 274
rect 17404 222 17410 274
rect 17534 222 17540 274
rect 17592 222 17598 274
rect 18016 150 18044 620
rect 18148 150 18176 620
rect 18376 500 18382 552
rect 18434 500 18440 552
rect 18612 274 18640 620
rect 18800 274 18828 620
rect 19000 376 19006 428
rect 19058 376 19064 428
rect 18594 222 18600 274
rect 18652 222 18658 274
rect 18782 222 18788 274
rect 18840 222 18846 274
rect 19264 150 19292 620
rect 19396 150 19424 620
rect 19624 500 19630 552
rect 19682 500 19688 552
rect 19860 274 19888 620
rect 20048 274 20076 620
rect 20248 376 20254 428
rect 20306 376 20312 428
rect 19842 222 19848 274
rect 19900 222 19906 274
rect 20030 222 20036 274
rect 20088 222 20094 274
rect 20512 150 20540 620
rect 20644 150 20672 620
rect 20872 500 20878 552
rect 20930 500 20936 552
rect 21108 274 21136 620
rect 21296 274 21324 620
rect 21496 376 21502 428
rect 21554 376 21560 428
rect 21090 222 21096 274
rect 21148 222 21154 274
rect 21278 222 21284 274
rect 21336 222 21342 274
rect 21760 150 21788 620
rect 21892 150 21920 620
rect 22120 500 22126 552
rect 22178 500 22184 552
rect 22356 274 22384 620
rect 22544 274 22572 620
rect 22744 376 22750 428
rect 22802 376 22808 428
rect 22338 222 22344 274
rect 22396 222 22402 274
rect 22526 222 22532 274
rect 22584 222 22590 274
rect 23008 150 23036 620
rect 23140 150 23168 620
rect 23368 500 23374 552
rect 23426 500 23432 552
rect 23604 274 23632 620
rect 23792 274 23820 620
rect 23992 376 23998 428
rect 24050 376 24056 428
rect 23586 222 23592 274
rect 23644 222 23650 274
rect 23774 222 23780 274
rect 23832 222 23838 274
rect 24256 150 24284 620
rect 24388 150 24416 620
rect 24616 500 24622 552
rect 24674 500 24680 552
rect 24852 274 24880 620
rect 25040 274 25068 620
rect 25240 376 25246 428
rect 25298 376 25304 428
rect 24834 222 24840 274
rect 24892 222 24898 274
rect 25022 222 25028 274
rect 25080 222 25086 274
rect 25504 150 25532 620
rect 25636 150 25664 620
rect 25864 500 25870 552
rect 25922 500 25928 552
rect 26100 274 26128 620
rect 26288 274 26316 620
rect 26488 376 26494 428
rect 26546 376 26552 428
rect 26082 222 26088 274
rect 26140 222 26146 274
rect 26270 222 26276 274
rect 26328 222 26334 274
rect 26752 150 26780 620
rect 26884 150 26912 620
rect 27112 500 27118 552
rect 27170 500 27176 552
rect 27348 274 27376 620
rect 27536 274 27564 620
rect 27736 376 27742 428
rect 27794 376 27800 428
rect 27330 222 27336 274
rect 27388 222 27394 274
rect 27518 222 27524 274
rect 27576 222 27582 274
rect 28000 150 28028 620
rect 28132 150 28160 620
rect 28360 500 28366 552
rect 28418 500 28424 552
rect 28596 274 28624 620
rect 28784 274 28812 620
rect 28984 376 28990 428
rect 29042 376 29048 428
rect 28578 222 28584 274
rect 28636 222 28642 274
rect 28766 222 28772 274
rect 28824 222 28830 274
rect 29248 150 29276 620
rect 29380 150 29408 620
rect 29608 500 29614 552
rect 29666 500 29672 552
rect 29844 274 29872 620
rect 30032 274 30060 620
rect 30232 376 30238 428
rect 30290 376 30296 428
rect 29826 222 29832 274
rect 29884 222 29890 274
rect 30014 222 30020 274
rect 30072 222 30078 274
rect 30496 150 30524 620
rect 30628 150 30656 620
rect 30856 500 30862 552
rect 30914 500 30920 552
rect 31092 274 31120 620
rect 31280 274 31308 620
rect 31480 376 31486 428
rect 31538 376 31544 428
rect 31074 222 31080 274
rect 31132 222 31138 274
rect 31262 222 31268 274
rect 31320 222 31326 274
rect 31744 150 31772 620
rect 31876 150 31904 620
rect 32104 500 32110 552
rect 32162 500 32168 552
rect 32340 274 32368 620
rect 32528 274 32556 620
rect 32728 376 32734 428
rect 32786 376 32792 428
rect 32322 222 32328 274
rect 32380 222 32386 274
rect 32510 222 32516 274
rect 32568 222 32574 274
rect 32992 150 33020 620
rect 33124 150 33152 620
rect 33352 500 33358 552
rect 33410 500 33416 552
rect 33588 274 33616 620
rect 33776 274 33804 620
rect 33976 376 33982 428
rect 34034 376 34040 428
rect 33570 222 33576 274
rect 33628 222 33634 274
rect 33758 222 33764 274
rect 33816 222 33822 274
rect 34240 150 34268 620
rect 34372 150 34400 620
rect 34600 500 34606 552
rect 34658 500 34664 552
rect 34836 274 34864 620
rect 35024 274 35052 620
rect 35224 376 35230 428
rect 35282 376 35288 428
rect 34818 222 34824 274
rect 34876 222 34882 274
rect 35006 222 35012 274
rect 35064 222 35070 274
rect 35488 150 35516 620
rect 35620 150 35648 620
rect 35848 500 35854 552
rect 35906 500 35912 552
rect 36084 274 36112 620
rect 36272 274 36300 620
rect 36472 376 36478 428
rect 36530 376 36536 428
rect 36066 222 36072 274
rect 36124 222 36130 274
rect 36254 222 36260 274
rect 36312 222 36318 274
rect 36736 150 36764 620
rect 36868 150 36896 620
rect 37096 500 37102 552
rect 37154 500 37160 552
rect 37332 274 37360 620
rect 37520 274 37548 620
rect 37720 376 37726 428
rect 37778 376 37784 428
rect 37314 222 37320 274
rect 37372 222 37378 274
rect 37502 222 37508 274
rect 37560 222 37566 274
rect 37984 150 38012 620
rect 38116 150 38144 620
rect 38344 500 38350 552
rect 38402 500 38408 552
rect 38580 274 38608 620
rect 38768 274 38796 620
rect 38968 376 38974 428
rect 39026 376 39032 428
rect 38562 222 38568 274
rect 38620 222 38626 274
rect 38750 222 38756 274
rect 38808 222 38814 274
rect 39232 150 39260 620
rect 39364 150 39392 620
rect 39592 500 39598 552
rect 39650 500 39656 552
rect 39828 274 39856 620
rect 39810 222 39816 274
rect 39868 222 39874 274
rect 526 98 532 150
rect 584 98 590 150
rect 658 98 664 150
rect 716 98 722 150
rect 1774 98 1780 150
rect 1832 98 1838 150
rect 1906 98 1912 150
rect 1964 98 1970 150
rect 3022 98 3028 150
rect 3080 98 3086 150
rect 3154 98 3160 150
rect 3212 98 3218 150
rect 4270 98 4276 150
rect 4328 98 4334 150
rect 4402 98 4408 150
rect 4460 98 4466 150
rect 5518 98 5524 150
rect 5576 98 5582 150
rect 5650 98 5656 150
rect 5708 98 5714 150
rect 6766 98 6772 150
rect 6824 98 6830 150
rect 6898 98 6904 150
rect 6956 98 6962 150
rect 8014 98 8020 150
rect 8072 98 8078 150
rect 8146 98 8152 150
rect 8204 98 8210 150
rect 9262 98 9268 150
rect 9320 98 9326 150
rect 9394 98 9400 150
rect 9452 98 9458 150
rect 10510 98 10516 150
rect 10568 98 10574 150
rect 10642 98 10648 150
rect 10700 98 10706 150
rect 11758 98 11764 150
rect 11816 98 11822 150
rect 11890 98 11896 150
rect 11948 98 11954 150
rect 13006 98 13012 150
rect 13064 98 13070 150
rect 13138 98 13144 150
rect 13196 98 13202 150
rect 14254 98 14260 150
rect 14312 98 14318 150
rect 14386 98 14392 150
rect 14444 98 14450 150
rect 15502 98 15508 150
rect 15560 98 15566 150
rect 15634 98 15640 150
rect 15692 98 15698 150
rect 16750 98 16756 150
rect 16808 98 16814 150
rect 16882 98 16888 150
rect 16940 98 16946 150
rect 17998 98 18004 150
rect 18056 98 18062 150
rect 18130 98 18136 150
rect 18188 98 18194 150
rect 19246 98 19252 150
rect 19304 98 19310 150
rect 19378 98 19384 150
rect 19436 98 19442 150
rect 20494 98 20500 150
rect 20552 98 20558 150
rect 20626 98 20632 150
rect 20684 98 20690 150
rect 21742 98 21748 150
rect 21800 98 21806 150
rect 21874 98 21880 150
rect 21932 98 21938 150
rect 22990 98 22996 150
rect 23048 98 23054 150
rect 23122 98 23128 150
rect 23180 98 23186 150
rect 24238 98 24244 150
rect 24296 98 24302 150
rect 24370 98 24376 150
rect 24428 98 24434 150
rect 25486 98 25492 150
rect 25544 98 25550 150
rect 25618 98 25624 150
rect 25676 98 25682 150
rect 26734 98 26740 150
rect 26792 98 26798 150
rect 26866 98 26872 150
rect 26924 98 26930 150
rect 27982 98 27988 150
rect 28040 98 28046 150
rect 28114 98 28120 150
rect 28172 98 28178 150
rect 29230 98 29236 150
rect 29288 98 29294 150
rect 29362 98 29368 150
rect 29420 98 29426 150
rect 30478 98 30484 150
rect 30536 98 30542 150
rect 30610 98 30616 150
rect 30668 98 30674 150
rect 31726 98 31732 150
rect 31784 98 31790 150
rect 31858 98 31864 150
rect 31916 98 31922 150
rect 32974 98 32980 150
rect 33032 98 33038 150
rect 33106 98 33112 150
rect 33164 98 33170 150
rect 34222 98 34228 150
rect 34280 98 34286 150
rect 34354 98 34360 150
rect 34412 98 34418 150
rect 35470 98 35476 150
rect 35528 98 35534 150
rect 35602 98 35608 150
rect 35660 98 35666 150
rect 36718 98 36724 150
rect 36776 98 36782 150
rect 36850 98 36856 150
rect 36908 98 36914 150
rect 37966 98 37972 150
rect 38024 98 38030 150
rect 38098 98 38104 150
rect 38156 98 38162 150
rect 39214 98 39220 150
rect 39272 98 39278 150
rect 39346 98 39352 150
rect 39404 98 39410 150
<< via1 >>
rect 286 419 338 428
rect 286 385 295 419
rect 295 385 329 419
rect 329 385 338 419
rect 286 376 338 385
rect 68 222 120 274
rect 910 543 962 552
rect 910 509 919 543
rect 919 509 953 543
rect 953 509 962 543
rect 910 500 962 509
rect 1534 419 1586 428
rect 1534 385 1543 419
rect 1543 385 1577 419
rect 1577 385 1586 419
rect 1534 376 1586 385
rect 1128 222 1180 274
rect 1316 222 1368 274
rect 2158 543 2210 552
rect 2158 509 2167 543
rect 2167 509 2201 543
rect 2201 509 2210 543
rect 2158 500 2210 509
rect 2782 419 2834 428
rect 2782 385 2791 419
rect 2791 385 2825 419
rect 2825 385 2834 419
rect 2782 376 2834 385
rect 2376 222 2428 274
rect 2564 222 2616 274
rect 3406 543 3458 552
rect 3406 509 3415 543
rect 3415 509 3449 543
rect 3449 509 3458 543
rect 3406 500 3458 509
rect 4030 419 4082 428
rect 4030 385 4039 419
rect 4039 385 4073 419
rect 4073 385 4082 419
rect 4030 376 4082 385
rect 3624 222 3676 274
rect 3812 222 3864 274
rect 4654 543 4706 552
rect 4654 509 4663 543
rect 4663 509 4697 543
rect 4697 509 4706 543
rect 4654 500 4706 509
rect 5278 419 5330 428
rect 5278 385 5287 419
rect 5287 385 5321 419
rect 5321 385 5330 419
rect 5278 376 5330 385
rect 4872 222 4924 274
rect 5060 222 5112 274
rect 5902 543 5954 552
rect 5902 509 5911 543
rect 5911 509 5945 543
rect 5945 509 5954 543
rect 5902 500 5954 509
rect 6526 419 6578 428
rect 6526 385 6535 419
rect 6535 385 6569 419
rect 6569 385 6578 419
rect 6526 376 6578 385
rect 6120 222 6172 274
rect 6308 222 6360 274
rect 7150 543 7202 552
rect 7150 509 7159 543
rect 7159 509 7193 543
rect 7193 509 7202 543
rect 7150 500 7202 509
rect 7774 419 7826 428
rect 7774 385 7783 419
rect 7783 385 7817 419
rect 7817 385 7826 419
rect 7774 376 7826 385
rect 7368 222 7420 274
rect 7556 222 7608 274
rect 8398 543 8450 552
rect 8398 509 8407 543
rect 8407 509 8441 543
rect 8441 509 8450 543
rect 8398 500 8450 509
rect 9022 419 9074 428
rect 9022 385 9031 419
rect 9031 385 9065 419
rect 9065 385 9074 419
rect 9022 376 9074 385
rect 8616 222 8668 274
rect 8804 222 8856 274
rect 9646 543 9698 552
rect 9646 509 9655 543
rect 9655 509 9689 543
rect 9689 509 9698 543
rect 9646 500 9698 509
rect 10270 419 10322 428
rect 10270 385 10279 419
rect 10279 385 10313 419
rect 10313 385 10322 419
rect 10270 376 10322 385
rect 9864 222 9916 274
rect 10052 222 10104 274
rect 10894 543 10946 552
rect 10894 509 10903 543
rect 10903 509 10937 543
rect 10937 509 10946 543
rect 10894 500 10946 509
rect 11518 419 11570 428
rect 11518 385 11527 419
rect 11527 385 11561 419
rect 11561 385 11570 419
rect 11518 376 11570 385
rect 11112 222 11164 274
rect 11300 222 11352 274
rect 12142 543 12194 552
rect 12142 509 12151 543
rect 12151 509 12185 543
rect 12185 509 12194 543
rect 12142 500 12194 509
rect 12766 419 12818 428
rect 12766 385 12775 419
rect 12775 385 12809 419
rect 12809 385 12818 419
rect 12766 376 12818 385
rect 12360 222 12412 274
rect 12548 222 12600 274
rect 13390 543 13442 552
rect 13390 509 13399 543
rect 13399 509 13433 543
rect 13433 509 13442 543
rect 13390 500 13442 509
rect 14014 419 14066 428
rect 14014 385 14023 419
rect 14023 385 14057 419
rect 14057 385 14066 419
rect 14014 376 14066 385
rect 13608 222 13660 274
rect 13796 222 13848 274
rect 14638 543 14690 552
rect 14638 509 14647 543
rect 14647 509 14681 543
rect 14681 509 14690 543
rect 14638 500 14690 509
rect 15262 419 15314 428
rect 15262 385 15271 419
rect 15271 385 15305 419
rect 15305 385 15314 419
rect 15262 376 15314 385
rect 14856 222 14908 274
rect 15044 222 15096 274
rect 15886 543 15938 552
rect 15886 509 15895 543
rect 15895 509 15929 543
rect 15929 509 15938 543
rect 15886 500 15938 509
rect 16510 419 16562 428
rect 16510 385 16519 419
rect 16519 385 16553 419
rect 16553 385 16562 419
rect 16510 376 16562 385
rect 16104 222 16156 274
rect 16292 222 16344 274
rect 17134 543 17186 552
rect 17134 509 17143 543
rect 17143 509 17177 543
rect 17177 509 17186 543
rect 17134 500 17186 509
rect 17758 419 17810 428
rect 17758 385 17767 419
rect 17767 385 17801 419
rect 17801 385 17810 419
rect 17758 376 17810 385
rect 17352 222 17404 274
rect 17540 222 17592 274
rect 18382 543 18434 552
rect 18382 509 18391 543
rect 18391 509 18425 543
rect 18425 509 18434 543
rect 18382 500 18434 509
rect 19006 419 19058 428
rect 19006 385 19015 419
rect 19015 385 19049 419
rect 19049 385 19058 419
rect 19006 376 19058 385
rect 18600 222 18652 274
rect 18788 222 18840 274
rect 19630 543 19682 552
rect 19630 509 19639 543
rect 19639 509 19673 543
rect 19673 509 19682 543
rect 19630 500 19682 509
rect 20254 419 20306 428
rect 20254 385 20263 419
rect 20263 385 20297 419
rect 20297 385 20306 419
rect 20254 376 20306 385
rect 19848 222 19900 274
rect 20036 222 20088 274
rect 20878 543 20930 552
rect 20878 509 20887 543
rect 20887 509 20921 543
rect 20921 509 20930 543
rect 20878 500 20930 509
rect 21502 419 21554 428
rect 21502 385 21511 419
rect 21511 385 21545 419
rect 21545 385 21554 419
rect 21502 376 21554 385
rect 21096 222 21148 274
rect 21284 222 21336 274
rect 22126 543 22178 552
rect 22126 509 22135 543
rect 22135 509 22169 543
rect 22169 509 22178 543
rect 22126 500 22178 509
rect 22750 419 22802 428
rect 22750 385 22759 419
rect 22759 385 22793 419
rect 22793 385 22802 419
rect 22750 376 22802 385
rect 22344 222 22396 274
rect 22532 222 22584 274
rect 23374 543 23426 552
rect 23374 509 23383 543
rect 23383 509 23417 543
rect 23417 509 23426 543
rect 23374 500 23426 509
rect 23998 419 24050 428
rect 23998 385 24007 419
rect 24007 385 24041 419
rect 24041 385 24050 419
rect 23998 376 24050 385
rect 23592 222 23644 274
rect 23780 222 23832 274
rect 24622 543 24674 552
rect 24622 509 24631 543
rect 24631 509 24665 543
rect 24665 509 24674 543
rect 24622 500 24674 509
rect 25246 419 25298 428
rect 25246 385 25255 419
rect 25255 385 25289 419
rect 25289 385 25298 419
rect 25246 376 25298 385
rect 24840 222 24892 274
rect 25028 222 25080 274
rect 25870 543 25922 552
rect 25870 509 25879 543
rect 25879 509 25913 543
rect 25913 509 25922 543
rect 25870 500 25922 509
rect 26494 419 26546 428
rect 26494 385 26503 419
rect 26503 385 26537 419
rect 26537 385 26546 419
rect 26494 376 26546 385
rect 26088 222 26140 274
rect 26276 222 26328 274
rect 27118 543 27170 552
rect 27118 509 27127 543
rect 27127 509 27161 543
rect 27161 509 27170 543
rect 27118 500 27170 509
rect 27742 419 27794 428
rect 27742 385 27751 419
rect 27751 385 27785 419
rect 27785 385 27794 419
rect 27742 376 27794 385
rect 27336 222 27388 274
rect 27524 222 27576 274
rect 28366 543 28418 552
rect 28366 509 28375 543
rect 28375 509 28409 543
rect 28409 509 28418 543
rect 28366 500 28418 509
rect 28990 419 29042 428
rect 28990 385 28999 419
rect 28999 385 29033 419
rect 29033 385 29042 419
rect 28990 376 29042 385
rect 28584 222 28636 274
rect 28772 222 28824 274
rect 29614 543 29666 552
rect 29614 509 29623 543
rect 29623 509 29657 543
rect 29657 509 29666 543
rect 29614 500 29666 509
rect 30238 419 30290 428
rect 30238 385 30247 419
rect 30247 385 30281 419
rect 30281 385 30290 419
rect 30238 376 30290 385
rect 29832 222 29884 274
rect 30020 222 30072 274
rect 30862 543 30914 552
rect 30862 509 30871 543
rect 30871 509 30905 543
rect 30905 509 30914 543
rect 30862 500 30914 509
rect 31486 419 31538 428
rect 31486 385 31495 419
rect 31495 385 31529 419
rect 31529 385 31538 419
rect 31486 376 31538 385
rect 31080 222 31132 274
rect 31268 222 31320 274
rect 32110 543 32162 552
rect 32110 509 32119 543
rect 32119 509 32153 543
rect 32153 509 32162 543
rect 32110 500 32162 509
rect 32734 419 32786 428
rect 32734 385 32743 419
rect 32743 385 32777 419
rect 32777 385 32786 419
rect 32734 376 32786 385
rect 32328 222 32380 274
rect 32516 222 32568 274
rect 33358 543 33410 552
rect 33358 509 33367 543
rect 33367 509 33401 543
rect 33401 509 33410 543
rect 33358 500 33410 509
rect 33982 419 34034 428
rect 33982 385 33991 419
rect 33991 385 34025 419
rect 34025 385 34034 419
rect 33982 376 34034 385
rect 33576 222 33628 274
rect 33764 222 33816 274
rect 34606 543 34658 552
rect 34606 509 34615 543
rect 34615 509 34649 543
rect 34649 509 34658 543
rect 34606 500 34658 509
rect 35230 419 35282 428
rect 35230 385 35239 419
rect 35239 385 35273 419
rect 35273 385 35282 419
rect 35230 376 35282 385
rect 34824 222 34876 274
rect 35012 222 35064 274
rect 35854 543 35906 552
rect 35854 509 35863 543
rect 35863 509 35897 543
rect 35897 509 35906 543
rect 35854 500 35906 509
rect 36478 419 36530 428
rect 36478 385 36487 419
rect 36487 385 36521 419
rect 36521 385 36530 419
rect 36478 376 36530 385
rect 36072 222 36124 274
rect 36260 222 36312 274
rect 37102 543 37154 552
rect 37102 509 37111 543
rect 37111 509 37145 543
rect 37145 509 37154 543
rect 37102 500 37154 509
rect 37726 419 37778 428
rect 37726 385 37735 419
rect 37735 385 37769 419
rect 37769 385 37778 419
rect 37726 376 37778 385
rect 37320 222 37372 274
rect 37508 222 37560 274
rect 38350 543 38402 552
rect 38350 509 38359 543
rect 38359 509 38393 543
rect 38393 509 38402 543
rect 38350 500 38402 509
rect 38974 419 39026 428
rect 38974 385 38983 419
rect 38983 385 39017 419
rect 39017 385 39026 419
rect 38974 376 39026 385
rect 38568 222 38620 274
rect 38756 222 38808 274
rect 39598 543 39650 552
rect 39598 509 39607 543
rect 39607 509 39641 543
rect 39641 509 39650 543
rect 39598 500 39650 509
rect 39816 222 39868 274
rect 532 98 584 150
rect 664 98 716 150
rect 1780 98 1832 150
rect 1912 98 1964 150
rect 3028 98 3080 150
rect 3160 98 3212 150
rect 4276 98 4328 150
rect 4408 98 4460 150
rect 5524 98 5576 150
rect 5656 98 5708 150
rect 6772 98 6824 150
rect 6904 98 6956 150
rect 8020 98 8072 150
rect 8152 98 8204 150
rect 9268 98 9320 150
rect 9400 98 9452 150
rect 10516 98 10568 150
rect 10648 98 10700 150
rect 11764 98 11816 150
rect 11896 98 11948 150
rect 13012 98 13064 150
rect 13144 98 13196 150
rect 14260 98 14312 150
rect 14392 98 14444 150
rect 15508 98 15560 150
rect 15640 98 15692 150
rect 16756 98 16808 150
rect 16888 98 16940 150
rect 18004 98 18056 150
rect 18136 98 18188 150
rect 19252 98 19304 150
rect 19384 98 19436 150
rect 20500 98 20552 150
rect 20632 98 20684 150
rect 21748 98 21800 150
rect 21880 98 21932 150
rect 22996 98 23048 150
rect 23128 98 23180 150
rect 24244 98 24296 150
rect 24376 98 24428 150
rect 25492 98 25544 150
rect 25624 98 25676 150
rect 26740 98 26792 150
rect 26872 98 26924 150
rect 27988 98 28040 150
rect 28120 98 28172 150
rect 29236 98 29288 150
rect 29368 98 29420 150
rect 30484 98 30536 150
rect 30616 98 30668 150
rect 31732 98 31784 150
rect 31864 98 31916 150
rect 32980 98 33032 150
rect 33112 98 33164 150
rect 34228 98 34280 150
rect 34360 98 34412 150
rect 35476 98 35528 150
rect 35608 98 35660 150
rect 36724 98 36776 150
rect 36856 98 36908 150
rect 37972 98 38024 150
rect 38104 98 38156 150
rect 39220 98 39272 150
rect 39352 98 39404 150
<< metal2 >>
rect 908 554 964 563
rect 908 489 964 498
rect 2156 554 2212 563
rect 2156 489 2212 498
rect 3404 554 3460 563
rect 3404 489 3460 498
rect 4652 554 4708 563
rect 4652 489 4708 498
rect 5900 554 5956 563
rect 5900 489 5956 498
rect 7148 554 7204 563
rect 7148 489 7204 498
rect 8396 554 8452 563
rect 8396 489 8452 498
rect 9644 554 9700 563
rect 9644 489 9700 498
rect 10892 554 10948 563
rect 10892 489 10948 498
rect 12140 554 12196 563
rect 12140 489 12196 498
rect 13388 554 13444 563
rect 13388 489 13444 498
rect 14636 554 14692 563
rect 14636 489 14692 498
rect 15884 554 15940 563
rect 15884 489 15940 498
rect 17132 554 17188 563
rect 17132 489 17188 498
rect 18380 554 18436 563
rect 18380 489 18436 498
rect 19628 554 19684 563
rect 19628 489 19684 498
rect 20876 554 20932 563
rect 20876 489 20932 498
rect 22124 554 22180 563
rect 22124 489 22180 498
rect 23372 554 23428 563
rect 23372 489 23428 498
rect 24620 554 24676 563
rect 24620 489 24676 498
rect 25868 554 25924 563
rect 25868 489 25924 498
rect 27116 554 27172 563
rect 27116 489 27172 498
rect 28364 554 28420 563
rect 28364 489 28420 498
rect 29612 554 29668 563
rect 29612 489 29668 498
rect 30860 554 30916 563
rect 30860 489 30916 498
rect 32108 554 32164 563
rect 32108 489 32164 498
rect 33356 554 33412 563
rect 33356 489 33412 498
rect 34604 554 34660 563
rect 34604 489 34660 498
rect 35852 554 35908 563
rect 35852 489 35908 498
rect 37100 554 37156 563
rect 37100 489 37156 498
rect 38348 554 38404 563
rect 38348 489 38404 498
rect 39596 554 39652 563
rect 39596 489 39652 498
rect 284 430 340 439
rect 284 365 340 374
rect 1532 430 1588 439
rect 1532 365 1588 374
rect 2780 430 2836 439
rect 2780 365 2836 374
rect 4028 430 4084 439
rect 4028 365 4084 374
rect 5276 430 5332 439
rect 5276 365 5332 374
rect 6524 430 6580 439
rect 6524 365 6580 374
rect 7772 430 7828 439
rect 7772 365 7828 374
rect 9020 430 9076 439
rect 9020 365 9076 374
rect 10268 430 10324 439
rect 10268 365 10324 374
rect 11516 430 11572 439
rect 11516 365 11572 374
rect 12764 430 12820 439
rect 12764 365 12820 374
rect 14012 430 14068 439
rect 14012 365 14068 374
rect 15260 430 15316 439
rect 15260 365 15316 374
rect 16508 430 16564 439
rect 16508 365 16564 374
rect 17756 430 17812 439
rect 17756 365 17812 374
rect 19004 430 19060 439
rect 19004 365 19060 374
rect 20252 430 20308 439
rect 20252 365 20308 374
rect 21500 430 21556 439
rect 21500 365 21556 374
rect 22748 430 22804 439
rect 22748 365 22804 374
rect 23996 430 24052 439
rect 23996 365 24052 374
rect 25244 430 25300 439
rect 25244 365 25300 374
rect 26492 430 26548 439
rect 26492 365 26548 374
rect 27740 430 27796 439
rect 27740 365 27796 374
rect 28988 430 29044 439
rect 28988 365 29044 374
rect 30236 430 30292 439
rect 30236 365 30292 374
rect 31484 430 31540 439
rect 31484 365 31540 374
rect 32732 430 32788 439
rect 32732 365 32788 374
rect 33980 430 34036 439
rect 33980 365 34036 374
rect 35228 430 35284 439
rect 35228 365 35284 374
rect 36476 430 36532 439
rect 36476 365 36532 374
rect 37724 430 37780 439
rect 37724 365 37780 374
rect 38972 430 39028 439
rect 38972 365 39028 374
rect 66 276 122 285
rect 66 211 122 220
rect 1126 276 1182 285
rect 1126 211 1182 220
rect 1314 276 1370 285
rect 1314 211 1370 220
rect 2374 276 2430 285
rect 2374 211 2430 220
rect 2562 276 2618 285
rect 2562 211 2618 220
rect 3622 276 3678 285
rect 3622 211 3678 220
rect 3810 276 3866 285
rect 3810 211 3866 220
rect 4870 276 4926 285
rect 4870 211 4926 220
rect 5058 276 5114 285
rect 5058 211 5114 220
rect 6118 276 6174 285
rect 6118 211 6174 220
rect 6306 276 6362 285
rect 6306 211 6362 220
rect 7366 276 7422 285
rect 7366 211 7422 220
rect 7554 276 7610 285
rect 7554 211 7610 220
rect 8614 276 8670 285
rect 8614 211 8670 220
rect 8802 276 8858 285
rect 8802 211 8858 220
rect 9862 276 9918 285
rect 9862 211 9918 220
rect 10050 276 10106 285
rect 10050 211 10106 220
rect 11110 276 11166 285
rect 11110 211 11166 220
rect 11298 276 11354 285
rect 11298 211 11354 220
rect 12358 276 12414 285
rect 12358 211 12414 220
rect 12546 276 12602 285
rect 12546 211 12602 220
rect 13606 276 13662 285
rect 13606 211 13662 220
rect 13794 276 13850 285
rect 13794 211 13850 220
rect 14854 276 14910 285
rect 14854 211 14910 220
rect 15042 276 15098 285
rect 15042 211 15098 220
rect 16102 276 16158 285
rect 16102 211 16158 220
rect 16290 276 16346 285
rect 16290 211 16346 220
rect 17350 276 17406 285
rect 17350 211 17406 220
rect 17538 276 17594 285
rect 17538 211 17594 220
rect 18598 276 18654 285
rect 18598 211 18654 220
rect 18786 276 18842 285
rect 18786 211 18842 220
rect 19846 276 19902 285
rect 19846 211 19902 220
rect 20034 276 20090 285
rect 20034 211 20090 220
rect 21094 276 21150 285
rect 21094 211 21150 220
rect 21282 276 21338 285
rect 21282 211 21338 220
rect 22342 276 22398 285
rect 22342 211 22398 220
rect 22530 276 22586 285
rect 22530 211 22586 220
rect 23590 276 23646 285
rect 23590 211 23646 220
rect 23778 276 23834 285
rect 23778 211 23834 220
rect 24838 276 24894 285
rect 24838 211 24894 220
rect 25026 276 25082 285
rect 25026 211 25082 220
rect 26086 276 26142 285
rect 26086 211 26142 220
rect 26274 276 26330 285
rect 26274 211 26330 220
rect 27334 276 27390 285
rect 27334 211 27390 220
rect 27522 276 27578 285
rect 27522 211 27578 220
rect 28582 276 28638 285
rect 28582 211 28638 220
rect 28770 276 28826 285
rect 28770 211 28826 220
rect 29830 276 29886 285
rect 29830 211 29886 220
rect 30018 276 30074 285
rect 30018 211 30074 220
rect 31078 276 31134 285
rect 31078 211 31134 220
rect 31266 276 31322 285
rect 31266 211 31322 220
rect 32326 276 32382 285
rect 32326 211 32382 220
rect 32514 276 32570 285
rect 32514 211 32570 220
rect 33574 276 33630 285
rect 33574 211 33630 220
rect 33762 276 33818 285
rect 33762 211 33818 220
rect 34822 276 34878 285
rect 34822 211 34878 220
rect 35010 276 35066 285
rect 35010 211 35066 220
rect 36070 276 36126 285
rect 36070 211 36126 220
rect 36258 276 36314 285
rect 36258 211 36314 220
rect 37318 276 37374 285
rect 37318 211 37374 220
rect 37506 276 37562 285
rect 37506 211 37562 220
rect 38566 276 38622 285
rect 38566 211 38622 220
rect 38754 276 38810 285
rect 38754 211 38810 220
rect 39814 276 39870 285
rect 39814 211 39870 220
rect 530 152 586 161
rect 530 87 586 96
rect 662 152 718 161
rect 662 87 718 96
rect 1778 152 1834 161
rect 1778 87 1834 96
rect 1910 152 1966 161
rect 1910 87 1966 96
rect 3026 152 3082 161
rect 3026 87 3082 96
rect 3158 152 3214 161
rect 3158 87 3214 96
rect 4274 152 4330 161
rect 4274 87 4330 96
rect 4406 152 4462 161
rect 4406 87 4462 96
rect 5522 152 5578 161
rect 5522 87 5578 96
rect 5654 152 5710 161
rect 5654 87 5710 96
rect 6770 152 6826 161
rect 6770 87 6826 96
rect 6902 152 6958 161
rect 6902 87 6958 96
rect 8018 152 8074 161
rect 8018 87 8074 96
rect 8150 152 8206 161
rect 8150 87 8206 96
rect 9266 152 9322 161
rect 9266 87 9322 96
rect 9398 152 9454 161
rect 9398 87 9454 96
rect 10514 152 10570 161
rect 10514 87 10570 96
rect 10646 152 10702 161
rect 10646 87 10702 96
rect 11762 152 11818 161
rect 11762 87 11818 96
rect 11894 152 11950 161
rect 11894 87 11950 96
rect 13010 152 13066 161
rect 13010 87 13066 96
rect 13142 152 13198 161
rect 13142 87 13198 96
rect 14258 152 14314 161
rect 14258 87 14314 96
rect 14390 152 14446 161
rect 14390 87 14446 96
rect 15506 152 15562 161
rect 15506 87 15562 96
rect 15638 152 15694 161
rect 15638 87 15694 96
rect 16754 152 16810 161
rect 16754 87 16810 96
rect 16886 152 16942 161
rect 16886 87 16942 96
rect 18002 152 18058 161
rect 18002 87 18058 96
rect 18134 152 18190 161
rect 18134 87 18190 96
rect 19250 152 19306 161
rect 19250 87 19306 96
rect 19382 152 19438 161
rect 19382 87 19438 96
rect 20498 152 20554 161
rect 20498 87 20554 96
rect 20630 152 20686 161
rect 20630 87 20686 96
rect 21746 152 21802 161
rect 21746 87 21802 96
rect 21878 152 21934 161
rect 21878 87 21934 96
rect 22994 152 23050 161
rect 22994 87 23050 96
rect 23126 152 23182 161
rect 23126 87 23182 96
rect 24242 152 24298 161
rect 24242 87 24298 96
rect 24374 152 24430 161
rect 24374 87 24430 96
rect 25490 152 25546 161
rect 25490 87 25546 96
rect 25622 152 25678 161
rect 25622 87 25678 96
rect 26738 152 26794 161
rect 26738 87 26794 96
rect 26870 152 26926 161
rect 26870 87 26926 96
rect 27986 152 28042 161
rect 27986 87 28042 96
rect 28118 152 28174 161
rect 28118 87 28174 96
rect 29234 152 29290 161
rect 29234 87 29290 96
rect 29366 152 29422 161
rect 29366 87 29422 96
rect 30482 152 30538 161
rect 30482 87 30538 96
rect 30614 152 30670 161
rect 30614 87 30670 96
rect 31730 152 31786 161
rect 31730 87 31786 96
rect 31862 152 31918 161
rect 31862 87 31918 96
rect 32978 152 33034 161
rect 32978 87 33034 96
rect 33110 152 33166 161
rect 33110 87 33166 96
rect 34226 152 34282 161
rect 34226 87 34282 96
rect 34358 152 34414 161
rect 34358 87 34414 96
rect 35474 152 35530 161
rect 35474 87 35530 96
rect 35606 152 35662 161
rect 35606 87 35662 96
rect 36722 152 36778 161
rect 36722 87 36778 96
rect 36854 152 36910 161
rect 36854 87 36910 96
rect 37970 152 38026 161
rect 37970 87 38026 96
rect 38102 152 38158 161
rect 38102 87 38158 96
rect 39218 152 39274 161
rect 39218 87 39274 96
rect 39350 152 39406 161
rect 39350 87 39406 96
<< via2 >>
rect 908 552 964 554
rect 908 500 910 552
rect 910 500 962 552
rect 962 500 964 552
rect 908 498 964 500
rect 2156 552 2212 554
rect 2156 500 2158 552
rect 2158 500 2210 552
rect 2210 500 2212 552
rect 2156 498 2212 500
rect 3404 552 3460 554
rect 3404 500 3406 552
rect 3406 500 3458 552
rect 3458 500 3460 552
rect 3404 498 3460 500
rect 4652 552 4708 554
rect 4652 500 4654 552
rect 4654 500 4706 552
rect 4706 500 4708 552
rect 4652 498 4708 500
rect 5900 552 5956 554
rect 5900 500 5902 552
rect 5902 500 5954 552
rect 5954 500 5956 552
rect 5900 498 5956 500
rect 7148 552 7204 554
rect 7148 500 7150 552
rect 7150 500 7202 552
rect 7202 500 7204 552
rect 7148 498 7204 500
rect 8396 552 8452 554
rect 8396 500 8398 552
rect 8398 500 8450 552
rect 8450 500 8452 552
rect 8396 498 8452 500
rect 9644 552 9700 554
rect 9644 500 9646 552
rect 9646 500 9698 552
rect 9698 500 9700 552
rect 9644 498 9700 500
rect 10892 552 10948 554
rect 10892 500 10894 552
rect 10894 500 10946 552
rect 10946 500 10948 552
rect 10892 498 10948 500
rect 12140 552 12196 554
rect 12140 500 12142 552
rect 12142 500 12194 552
rect 12194 500 12196 552
rect 12140 498 12196 500
rect 13388 552 13444 554
rect 13388 500 13390 552
rect 13390 500 13442 552
rect 13442 500 13444 552
rect 13388 498 13444 500
rect 14636 552 14692 554
rect 14636 500 14638 552
rect 14638 500 14690 552
rect 14690 500 14692 552
rect 14636 498 14692 500
rect 15884 552 15940 554
rect 15884 500 15886 552
rect 15886 500 15938 552
rect 15938 500 15940 552
rect 15884 498 15940 500
rect 17132 552 17188 554
rect 17132 500 17134 552
rect 17134 500 17186 552
rect 17186 500 17188 552
rect 17132 498 17188 500
rect 18380 552 18436 554
rect 18380 500 18382 552
rect 18382 500 18434 552
rect 18434 500 18436 552
rect 18380 498 18436 500
rect 19628 552 19684 554
rect 19628 500 19630 552
rect 19630 500 19682 552
rect 19682 500 19684 552
rect 19628 498 19684 500
rect 20876 552 20932 554
rect 20876 500 20878 552
rect 20878 500 20930 552
rect 20930 500 20932 552
rect 20876 498 20932 500
rect 22124 552 22180 554
rect 22124 500 22126 552
rect 22126 500 22178 552
rect 22178 500 22180 552
rect 22124 498 22180 500
rect 23372 552 23428 554
rect 23372 500 23374 552
rect 23374 500 23426 552
rect 23426 500 23428 552
rect 23372 498 23428 500
rect 24620 552 24676 554
rect 24620 500 24622 552
rect 24622 500 24674 552
rect 24674 500 24676 552
rect 24620 498 24676 500
rect 25868 552 25924 554
rect 25868 500 25870 552
rect 25870 500 25922 552
rect 25922 500 25924 552
rect 25868 498 25924 500
rect 27116 552 27172 554
rect 27116 500 27118 552
rect 27118 500 27170 552
rect 27170 500 27172 552
rect 27116 498 27172 500
rect 28364 552 28420 554
rect 28364 500 28366 552
rect 28366 500 28418 552
rect 28418 500 28420 552
rect 28364 498 28420 500
rect 29612 552 29668 554
rect 29612 500 29614 552
rect 29614 500 29666 552
rect 29666 500 29668 552
rect 29612 498 29668 500
rect 30860 552 30916 554
rect 30860 500 30862 552
rect 30862 500 30914 552
rect 30914 500 30916 552
rect 30860 498 30916 500
rect 32108 552 32164 554
rect 32108 500 32110 552
rect 32110 500 32162 552
rect 32162 500 32164 552
rect 32108 498 32164 500
rect 33356 552 33412 554
rect 33356 500 33358 552
rect 33358 500 33410 552
rect 33410 500 33412 552
rect 33356 498 33412 500
rect 34604 552 34660 554
rect 34604 500 34606 552
rect 34606 500 34658 552
rect 34658 500 34660 552
rect 34604 498 34660 500
rect 35852 552 35908 554
rect 35852 500 35854 552
rect 35854 500 35906 552
rect 35906 500 35908 552
rect 35852 498 35908 500
rect 37100 552 37156 554
rect 37100 500 37102 552
rect 37102 500 37154 552
rect 37154 500 37156 552
rect 37100 498 37156 500
rect 38348 552 38404 554
rect 38348 500 38350 552
rect 38350 500 38402 552
rect 38402 500 38404 552
rect 38348 498 38404 500
rect 39596 552 39652 554
rect 39596 500 39598 552
rect 39598 500 39650 552
rect 39650 500 39652 552
rect 39596 498 39652 500
rect 284 428 340 430
rect 284 376 286 428
rect 286 376 338 428
rect 338 376 340 428
rect 284 374 340 376
rect 1532 428 1588 430
rect 1532 376 1534 428
rect 1534 376 1586 428
rect 1586 376 1588 428
rect 1532 374 1588 376
rect 2780 428 2836 430
rect 2780 376 2782 428
rect 2782 376 2834 428
rect 2834 376 2836 428
rect 2780 374 2836 376
rect 4028 428 4084 430
rect 4028 376 4030 428
rect 4030 376 4082 428
rect 4082 376 4084 428
rect 4028 374 4084 376
rect 5276 428 5332 430
rect 5276 376 5278 428
rect 5278 376 5330 428
rect 5330 376 5332 428
rect 5276 374 5332 376
rect 6524 428 6580 430
rect 6524 376 6526 428
rect 6526 376 6578 428
rect 6578 376 6580 428
rect 6524 374 6580 376
rect 7772 428 7828 430
rect 7772 376 7774 428
rect 7774 376 7826 428
rect 7826 376 7828 428
rect 7772 374 7828 376
rect 9020 428 9076 430
rect 9020 376 9022 428
rect 9022 376 9074 428
rect 9074 376 9076 428
rect 9020 374 9076 376
rect 10268 428 10324 430
rect 10268 376 10270 428
rect 10270 376 10322 428
rect 10322 376 10324 428
rect 10268 374 10324 376
rect 11516 428 11572 430
rect 11516 376 11518 428
rect 11518 376 11570 428
rect 11570 376 11572 428
rect 11516 374 11572 376
rect 12764 428 12820 430
rect 12764 376 12766 428
rect 12766 376 12818 428
rect 12818 376 12820 428
rect 12764 374 12820 376
rect 14012 428 14068 430
rect 14012 376 14014 428
rect 14014 376 14066 428
rect 14066 376 14068 428
rect 14012 374 14068 376
rect 15260 428 15316 430
rect 15260 376 15262 428
rect 15262 376 15314 428
rect 15314 376 15316 428
rect 15260 374 15316 376
rect 16508 428 16564 430
rect 16508 376 16510 428
rect 16510 376 16562 428
rect 16562 376 16564 428
rect 16508 374 16564 376
rect 17756 428 17812 430
rect 17756 376 17758 428
rect 17758 376 17810 428
rect 17810 376 17812 428
rect 17756 374 17812 376
rect 19004 428 19060 430
rect 19004 376 19006 428
rect 19006 376 19058 428
rect 19058 376 19060 428
rect 19004 374 19060 376
rect 20252 428 20308 430
rect 20252 376 20254 428
rect 20254 376 20306 428
rect 20306 376 20308 428
rect 20252 374 20308 376
rect 21500 428 21556 430
rect 21500 376 21502 428
rect 21502 376 21554 428
rect 21554 376 21556 428
rect 21500 374 21556 376
rect 22748 428 22804 430
rect 22748 376 22750 428
rect 22750 376 22802 428
rect 22802 376 22804 428
rect 22748 374 22804 376
rect 23996 428 24052 430
rect 23996 376 23998 428
rect 23998 376 24050 428
rect 24050 376 24052 428
rect 23996 374 24052 376
rect 25244 428 25300 430
rect 25244 376 25246 428
rect 25246 376 25298 428
rect 25298 376 25300 428
rect 25244 374 25300 376
rect 26492 428 26548 430
rect 26492 376 26494 428
rect 26494 376 26546 428
rect 26546 376 26548 428
rect 26492 374 26548 376
rect 27740 428 27796 430
rect 27740 376 27742 428
rect 27742 376 27794 428
rect 27794 376 27796 428
rect 27740 374 27796 376
rect 28988 428 29044 430
rect 28988 376 28990 428
rect 28990 376 29042 428
rect 29042 376 29044 428
rect 28988 374 29044 376
rect 30236 428 30292 430
rect 30236 376 30238 428
rect 30238 376 30290 428
rect 30290 376 30292 428
rect 30236 374 30292 376
rect 31484 428 31540 430
rect 31484 376 31486 428
rect 31486 376 31538 428
rect 31538 376 31540 428
rect 31484 374 31540 376
rect 32732 428 32788 430
rect 32732 376 32734 428
rect 32734 376 32786 428
rect 32786 376 32788 428
rect 32732 374 32788 376
rect 33980 428 34036 430
rect 33980 376 33982 428
rect 33982 376 34034 428
rect 34034 376 34036 428
rect 33980 374 34036 376
rect 35228 428 35284 430
rect 35228 376 35230 428
rect 35230 376 35282 428
rect 35282 376 35284 428
rect 35228 374 35284 376
rect 36476 428 36532 430
rect 36476 376 36478 428
rect 36478 376 36530 428
rect 36530 376 36532 428
rect 36476 374 36532 376
rect 37724 428 37780 430
rect 37724 376 37726 428
rect 37726 376 37778 428
rect 37778 376 37780 428
rect 37724 374 37780 376
rect 38972 428 39028 430
rect 38972 376 38974 428
rect 38974 376 39026 428
rect 39026 376 39028 428
rect 38972 374 39028 376
rect 66 274 122 276
rect 66 222 68 274
rect 68 222 120 274
rect 120 222 122 274
rect 66 220 122 222
rect 1126 274 1182 276
rect 1126 222 1128 274
rect 1128 222 1180 274
rect 1180 222 1182 274
rect 1126 220 1182 222
rect 1314 274 1370 276
rect 1314 222 1316 274
rect 1316 222 1368 274
rect 1368 222 1370 274
rect 1314 220 1370 222
rect 2374 274 2430 276
rect 2374 222 2376 274
rect 2376 222 2428 274
rect 2428 222 2430 274
rect 2374 220 2430 222
rect 2562 274 2618 276
rect 2562 222 2564 274
rect 2564 222 2616 274
rect 2616 222 2618 274
rect 2562 220 2618 222
rect 3622 274 3678 276
rect 3622 222 3624 274
rect 3624 222 3676 274
rect 3676 222 3678 274
rect 3622 220 3678 222
rect 3810 274 3866 276
rect 3810 222 3812 274
rect 3812 222 3864 274
rect 3864 222 3866 274
rect 3810 220 3866 222
rect 4870 274 4926 276
rect 4870 222 4872 274
rect 4872 222 4924 274
rect 4924 222 4926 274
rect 4870 220 4926 222
rect 5058 274 5114 276
rect 5058 222 5060 274
rect 5060 222 5112 274
rect 5112 222 5114 274
rect 5058 220 5114 222
rect 6118 274 6174 276
rect 6118 222 6120 274
rect 6120 222 6172 274
rect 6172 222 6174 274
rect 6118 220 6174 222
rect 6306 274 6362 276
rect 6306 222 6308 274
rect 6308 222 6360 274
rect 6360 222 6362 274
rect 6306 220 6362 222
rect 7366 274 7422 276
rect 7366 222 7368 274
rect 7368 222 7420 274
rect 7420 222 7422 274
rect 7366 220 7422 222
rect 7554 274 7610 276
rect 7554 222 7556 274
rect 7556 222 7608 274
rect 7608 222 7610 274
rect 7554 220 7610 222
rect 8614 274 8670 276
rect 8614 222 8616 274
rect 8616 222 8668 274
rect 8668 222 8670 274
rect 8614 220 8670 222
rect 8802 274 8858 276
rect 8802 222 8804 274
rect 8804 222 8856 274
rect 8856 222 8858 274
rect 8802 220 8858 222
rect 9862 274 9918 276
rect 9862 222 9864 274
rect 9864 222 9916 274
rect 9916 222 9918 274
rect 9862 220 9918 222
rect 10050 274 10106 276
rect 10050 222 10052 274
rect 10052 222 10104 274
rect 10104 222 10106 274
rect 10050 220 10106 222
rect 11110 274 11166 276
rect 11110 222 11112 274
rect 11112 222 11164 274
rect 11164 222 11166 274
rect 11110 220 11166 222
rect 11298 274 11354 276
rect 11298 222 11300 274
rect 11300 222 11352 274
rect 11352 222 11354 274
rect 11298 220 11354 222
rect 12358 274 12414 276
rect 12358 222 12360 274
rect 12360 222 12412 274
rect 12412 222 12414 274
rect 12358 220 12414 222
rect 12546 274 12602 276
rect 12546 222 12548 274
rect 12548 222 12600 274
rect 12600 222 12602 274
rect 12546 220 12602 222
rect 13606 274 13662 276
rect 13606 222 13608 274
rect 13608 222 13660 274
rect 13660 222 13662 274
rect 13606 220 13662 222
rect 13794 274 13850 276
rect 13794 222 13796 274
rect 13796 222 13848 274
rect 13848 222 13850 274
rect 13794 220 13850 222
rect 14854 274 14910 276
rect 14854 222 14856 274
rect 14856 222 14908 274
rect 14908 222 14910 274
rect 14854 220 14910 222
rect 15042 274 15098 276
rect 15042 222 15044 274
rect 15044 222 15096 274
rect 15096 222 15098 274
rect 15042 220 15098 222
rect 16102 274 16158 276
rect 16102 222 16104 274
rect 16104 222 16156 274
rect 16156 222 16158 274
rect 16102 220 16158 222
rect 16290 274 16346 276
rect 16290 222 16292 274
rect 16292 222 16344 274
rect 16344 222 16346 274
rect 16290 220 16346 222
rect 17350 274 17406 276
rect 17350 222 17352 274
rect 17352 222 17404 274
rect 17404 222 17406 274
rect 17350 220 17406 222
rect 17538 274 17594 276
rect 17538 222 17540 274
rect 17540 222 17592 274
rect 17592 222 17594 274
rect 17538 220 17594 222
rect 18598 274 18654 276
rect 18598 222 18600 274
rect 18600 222 18652 274
rect 18652 222 18654 274
rect 18598 220 18654 222
rect 18786 274 18842 276
rect 18786 222 18788 274
rect 18788 222 18840 274
rect 18840 222 18842 274
rect 18786 220 18842 222
rect 19846 274 19902 276
rect 19846 222 19848 274
rect 19848 222 19900 274
rect 19900 222 19902 274
rect 19846 220 19902 222
rect 20034 274 20090 276
rect 20034 222 20036 274
rect 20036 222 20088 274
rect 20088 222 20090 274
rect 20034 220 20090 222
rect 21094 274 21150 276
rect 21094 222 21096 274
rect 21096 222 21148 274
rect 21148 222 21150 274
rect 21094 220 21150 222
rect 21282 274 21338 276
rect 21282 222 21284 274
rect 21284 222 21336 274
rect 21336 222 21338 274
rect 21282 220 21338 222
rect 22342 274 22398 276
rect 22342 222 22344 274
rect 22344 222 22396 274
rect 22396 222 22398 274
rect 22342 220 22398 222
rect 22530 274 22586 276
rect 22530 222 22532 274
rect 22532 222 22584 274
rect 22584 222 22586 274
rect 22530 220 22586 222
rect 23590 274 23646 276
rect 23590 222 23592 274
rect 23592 222 23644 274
rect 23644 222 23646 274
rect 23590 220 23646 222
rect 23778 274 23834 276
rect 23778 222 23780 274
rect 23780 222 23832 274
rect 23832 222 23834 274
rect 23778 220 23834 222
rect 24838 274 24894 276
rect 24838 222 24840 274
rect 24840 222 24892 274
rect 24892 222 24894 274
rect 24838 220 24894 222
rect 25026 274 25082 276
rect 25026 222 25028 274
rect 25028 222 25080 274
rect 25080 222 25082 274
rect 25026 220 25082 222
rect 26086 274 26142 276
rect 26086 222 26088 274
rect 26088 222 26140 274
rect 26140 222 26142 274
rect 26086 220 26142 222
rect 26274 274 26330 276
rect 26274 222 26276 274
rect 26276 222 26328 274
rect 26328 222 26330 274
rect 26274 220 26330 222
rect 27334 274 27390 276
rect 27334 222 27336 274
rect 27336 222 27388 274
rect 27388 222 27390 274
rect 27334 220 27390 222
rect 27522 274 27578 276
rect 27522 222 27524 274
rect 27524 222 27576 274
rect 27576 222 27578 274
rect 27522 220 27578 222
rect 28582 274 28638 276
rect 28582 222 28584 274
rect 28584 222 28636 274
rect 28636 222 28638 274
rect 28582 220 28638 222
rect 28770 274 28826 276
rect 28770 222 28772 274
rect 28772 222 28824 274
rect 28824 222 28826 274
rect 28770 220 28826 222
rect 29830 274 29886 276
rect 29830 222 29832 274
rect 29832 222 29884 274
rect 29884 222 29886 274
rect 29830 220 29886 222
rect 30018 274 30074 276
rect 30018 222 30020 274
rect 30020 222 30072 274
rect 30072 222 30074 274
rect 30018 220 30074 222
rect 31078 274 31134 276
rect 31078 222 31080 274
rect 31080 222 31132 274
rect 31132 222 31134 274
rect 31078 220 31134 222
rect 31266 274 31322 276
rect 31266 222 31268 274
rect 31268 222 31320 274
rect 31320 222 31322 274
rect 31266 220 31322 222
rect 32326 274 32382 276
rect 32326 222 32328 274
rect 32328 222 32380 274
rect 32380 222 32382 274
rect 32326 220 32382 222
rect 32514 274 32570 276
rect 32514 222 32516 274
rect 32516 222 32568 274
rect 32568 222 32570 274
rect 32514 220 32570 222
rect 33574 274 33630 276
rect 33574 222 33576 274
rect 33576 222 33628 274
rect 33628 222 33630 274
rect 33574 220 33630 222
rect 33762 274 33818 276
rect 33762 222 33764 274
rect 33764 222 33816 274
rect 33816 222 33818 274
rect 33762 220 33818 222
rect 34822 274 34878 276
rect 34822 222 34824 274
rect 34824 222 34876 274
rect 34876 222 34878 274
rect 34822 220 34878 222
rect 35010 274 35066 276
rect 35010 222 35012 274
rect 35012 222 35064 274
rect 35064 222 35066 274
rect 35010 220 35066 222
rect 36070 274 36126 276
rect 36070 222 36072 274
rect 36072 222 36124 274
rect 36124 222 36126 274
rect 36070 220 36126 222
rect 36258 274 36314 276
rect 36258 222 36260 274
rect 36260 222 36312 274
rect 36312 222 36314 274
rect 36258 220 36314 222
rect 37318 274 37374 276
rect 37318 222 37320 274
rect 37320 222 37372 274
rect 37372 222 37374 274
rect 37318 220 37374 222
rect 37506 274 37562 276
rect 37506 222 37508 274
rect 37508 222 37560 274
rect 37560 222 37562 274
rect 37506 220 37562 222
rect 38566 274 38622 276
rect 38566 222 38568 274
rect 38568 222 38620 274
rect 38620 222 38622 274
rect 38566 220 38622 222
rect 38754 274 38810 276
rect 38754 222 38756 274
rect 38756 222 38808 274
rect 38808 222 38810 274
rect 38754 220 38810 222
rect 39814 274 39870 276
rect 39814 222 39816 274
rect 39816 222 39868 274
rect 39868 222 39870 274
rect 39814 220 39870 222
rect 530 150 586 152
rect 530 98 532 150
rect 532 98 584 150
rect 584 98 586 150
rect 530 96 586 98
rect 662 150 718 152
rect 662 98 664 150
rect 664 98 716 150
rect 716 98 718 150
rect 662 96 718 98
rect 1778 150 1834 152
rect 1778 98 1780 150
rect 1780 98 1832 150
rect 1832 98 1834 150
rect 1778 96 1834 98
rect 1910 150 1966 152
rect 1910 98 1912 150
rect 1912 98 1964 150
rect 1964 98 1966 150
rect 1910 96 1966 98
rect 3026 150 3082 152
rect 3026 98 3028 150
rect 3028 98 3080 150
rect 3080 98 3082 150
rect 3026 96 3082 98
rect 3158 150 3214 152
rect 3158 98 3160 150
rect 3160 98 3212 150
rect 3212 98 3214 150
rect 3158 96 3214 98
rect 4274 150 4330 152
rect 4274 98 4276 150
rect 4276 98 4328 150
rect 4328 98 4330 150
rect 4274 96 4330 98
rect 4406 150 4462 152
rect 4406 98 4408 150
rect 4408 98 4460 150
rect 4460 98 4462 150
rect 4406 96 4462 98
rect 5522 150 5578 152
rect 5522 98 5524 150
rect 5524 98 5576 150
rect 5576 98 5578 150
rect 5522 96 5578 98
rect 5654 150 5710 152
rect 5654 98 5656 150
rect 5656 98 5708 150
rect 5708 98 5710 150
rect 5654 96 5710 98
rect 6770 150 6826 152
rect 6770 98 6772 150
rect 6772 98 6824 150
rect 6824 98 6826 150
rect 6770 96 6826 98
rect 6902 150 6958 152
rect 6902 98 6904 150
rect 6904 98 6956 150
rect 6956 98 6958 150
rect 6902 96 6958 98
rect 8018 150 8074 152
rect 8018 98 8020 150
rect 8020 98 8072 150
rect 8072 98 8074 150
rect 8018 96 8074 98
rect 8150 150 8206 152
rect 8150 98 8152 150
rect 8152 98 8204 150
rect 8204 98 8206 150
rect 8150 96 8206 98
rect 9266 150 9322 152
rect 9266 98 9268 150
rect 9268 98 9320 150
rect 9320 98 9322 150
rect 9266 96 9322 98
rect 9398 150 9454 152
rect 9398 98 9400 150
rect 9400 98 9452 150
rect 9452 98 9454 150
rect 9398 96 9454 98
rect 10514 150 10570 152
rect 10514 98 10516 150
rect 10516 98 10568 150
rect 10568 98 10570 150
rect 10514 96 10570 98
rect 10646 150 10702 152
rect 10646 98 10648 150
rect 10648 98 10700 150
rect 10700 98 10702 150
rect 10646 96 10702 98
rect 11762 150 11818 152
rect 11762 98 11764 150
rect 11764 98 11816 150
rect 11816 98 11818 150
rect 11762 96 11818 98
rect 11894 150 11950 152
rect 11894 98 11896 150
rect 11896 98 11948 150
rect 11948 98 11950 150
rect 11894 96 11950 98
rect 13010 150 13066 152
rect 13010 98 13012 150
rect 13012 98 13064 150
rect 13064 98 13066 150
rect 13010 96 13066 98
rect 13142 150 13198 152
rect 13142 98 13144 150
rect 13144 98 13196 150
rect 13196 98 13198 150
rect 13142 96 13198 98
rect 14258 150 14314 152
rect 14258 98 14260 150
rect 14260 98 14312 150
rect 14312 98 14314 150
rect 14258 96 14314 98
rect 14390 150 14446 152
rect 14390 98 14392 150
rect 14392 98 14444 150
rect 14444 98 14446 150
rect 14390 96 14446 98
rect 15506 150 15562 152
rect 15506 98 15508 150
rect 15508 98 15560 150
rect 15560 98 15562 150
rect 15506 96 15562 98
rect 15638 150 15694 152
rect 15638 98 15640 150
rect 15640 98 15692 150
rect 15692 98 15694 150
rect 15638 96 15694 98
rect 16754 150 16810 152
rect 16754 98 16756 150
rect 16756 98 16808 150
rect 16808 98 16810 150
rect 16754 96 16810 98
rect 16886 150 16942 152
rect 16886 98 16888 150
rect 16888 98 16940 150
rect 16940 98 16942 150
rect 16886 96 16942 98
rect 18002 150 18058 152
rect 18002 98 18004 150
rect 18004 98 18056 150
rect 18056 98 18058 150
rect 18002 96 18058 98
rect 18134 150 18190 152
rect 18134 98 18136 150
rect 18136 98 18188 150
rect 18188 98 18190 150
rect 18134 96 18190 98
rect 19250 150 19306 152
rect 19250 98 19252 150
rect 19252 98 19304 150
rect 19304 98 19306 150
rect 19250 96 19306 98
rect 19382 150 19438 152
rect 19382 98 19384 150
rect 19384 98 19436 150
rect 19436 98 19438 150
rect 19382 96 19438 98
rect 20498 150 20554 152
rect 20498 98 20500 150
rect 20500 98 20552 150
rect 20552 98 20554 150
rect 20498 96 20554 98
rect 20630 150 20686 152
rect 20630 98 20632 150
rect 20632 98 20684 150
rect 20684 98 20686 150
rect 20630 96 20686 98
rect 21746 150 21802 152
rect 21746 98 21748 150
rect 21748 98 21800 150
rect 21800 98 21802 150
rect 21746 96 21802 98
rect 21878 150 21934 152
rect 21878 98 21880 150
rect 21880 98 21932 150
rect 21932 98 21934 150
rect 21878 96 21934 98
rect 22994 150 23050 152
rect 22994 98 22996 150
rect 22996 98 23048 150
rect 23048 98 23050 150
rect 22994 96 23050 98
rect 23126 150 23182 152
rect 23126 98 23128 150
rect 23128 98 23180 150
rect 23180 98 23182 150
rect 23126 96 23182 98
rect 24242 150 24298 152
rect 24242 98 24244 150
rect 24244 98 24296 150
rect 24296 98 24298 150
rect 24242 96 24298 98
rect 24374 150 24430 152
rect 24374 98 24376 150
rect 24376 98 24428 150
rect 24428 98 24430 150
rect 24374 96 24430 98
rect 25490 150 25546 152
rect 25490 98 25492 150
rect 25492 98 25544 150
rect 25544 98 25546 150
rect 25490 96 25546 98
rect 25622 150 25678 152
rect 25622 98 25624 150
rect 25624 98 25676 150
rect 25676 98 25678 150
rect 25622 96 25678 98
rect 26738 150 26794 152
rect 26738 98 26740 150
rect 26740 98 26792 150
rect 26792 98 26794 150
rect 26738 96 26794 98
rect 26870 150 26926 152
rect 26870 98 26872 150
rect 26872 98 26924 150
rect 26924 98 26926 150
rect 26870 96 26926 98
rect 27986 150 28042 152
rect 27986 98 27988 150
rect 27988 98 28040 150
rect 28040 98 28042 150
rect 27986 96 28042 98
rect 28118 150 28174 152
rect 28118 98 28120 150
rect 28120 98 28172 150
rect 28172 98 28174 150
rect 28118 96 28174 98
rect 29234 150 29290 152
rect 29234 98 29236 150
rect 29236 98 29288 150
rect 29288 98 29290 150
rect 29234 96 29290 98
rect 29366 150 29422 152
rect 29366 98 29368 150
rect 29368 98 29420 150
rect 29420 98 29422 150
rect 29366 96 29422 98
rect 30482 150 30538 152
rect 30482 98 30484 150
rect 30484 98 30536 150
rect 30536 98 30538 150
rect 30482 96 30538 98
rect 30614 150 30670 152
rect 30614 98 30616 150
rect 30616 98 30668 150
rect 30668 98 30670 150
rect 30614 96 30670 98
rect 31730 150 31786 152
rect 31730 98 31732 150
rect 31732 98 31784 150
rect 31784 98 31786 150
rect 31730 96 31786 98
rect 31862 150 31918 152
rect 31862 98 31864 150
rect 31864 98 31916 150
rect 31916 98 31918 150
rect 31862 96 31918 98
rect 32978 150 33034 152
rect 32978 98 32980 150
rect 32980 98 33032 150
rect 33032 98 33034 150
rect 32978 96 33034 98
rect 33110 150 33166 152
rect 33110 98 33112 150
rect 33112 98 33164 150
rect 33164 98 33166 150
rect 33110 96 33166 98
rect 34226 150 34282 152
rect 34226 98 34228 150
rect 34228 98 34280 150
rect 34280 98 34282 150
rect 34226 96 34282 98
rect 34358 150 34414 152
rect 34358 98 34360 150
rect 34360 98 34412 150
rect 34412 98 34414 150
rect 34358 96 34414 98
rect 35474 150 35530 152
rect 35474 98 35476 150
rect 35476 98 35528 150
rect 35528 98 35530 150
rect 35474 96 35530 98
rect 35606 150 35662 152
rect 35606 98 35608 150
rect 35608 98 35660 150
rect 35660 98 35662 150
rect 35606 96 35662 98
rect 36722 150 36778 152
rect 36722 98 36724 150
rect 36724 98 36776 150
rect 36776 98 36778 150
rect 36722 96 36778 98
rect 36854 150 36910 152
rect 36854 98 36856 150
rect 36856 98 36908 150
rect 36908 98 36910 150
rect 36854 96 36910 98
rect 37970 150 38026 152
rect 37970 98 37972 150
rect 37972 98 38024 150
rect 38024 98 38026 150
rect 37970 96 38026 98
rect 38102 150 38158 152
rect 38102 98 38104 150
rect 38104 98 38156 150
rect 38156 98 38158 150
rect 38102 96 38158 98
rect 39218 150 39274 152
rect 39218 98 39220 150
rect 39220 98 39272 150
rect 39272 98 39274 150
rect 39218 96 39274 98
rect 39350 150 39406 152
rect 39350 98 39352 150
rect 39352 98 39404 150
rect 39404 98 39406 150
rect 39350 96 39406 98
<< metal3 >>
rect 575 1258 673 1356
rect 1823 1258 1921 1356
rect 3071 1258 3169 1356
rect 4319 1258 4417 1356
rect 5567 1258 5665 1356
rect 6815 1258 6913 1356
rect 8063 1258 8161 1356
rect 9311 1258 9409 1356
rect 10559 1258 10657 1356
rect 11807 1258 11905 1356
rect 13055 1258 13153 1356
rect 14303 1258 14401 1356
rect 15551 1258 15649 1356
rect 16799 1258 16897 1356
rect 18047 1258 18145 1356
rect 19295 1258 19393 1356
rect 20543 1258 20641 1356
rect 21791 1258 21889 1356
rect 23039 1258 23137 1356
rect 24287 1258 24385 1356
rect 25535 1258 25633 1356
rect 26783 1258 26881 1356
rect 28031 1258 28129 1356
rect 29279 1258 29377 1356
rect 30527 1258 30625 1356
rect 31775 1258 31873 1356
rect 33023 1258 33121 1356
rect 34271 1258 34369 1356
rect 35519 1258 35617 1356
rect 36767 1258 36865 1356
rect 38015 1258 38113 1356
rect 39263 1258 39361 1356
rect 903 556 969 559
rect 2151 556 2217 559
rect 3399 556 3465 559
rect 4647 556 4713 559
rect 5895 556 5961 559
rect 7143 556 7209 559
rect 8391 556 8457 559
rect 9639 556 9705 559
rect 10887 556 10953 559
rect 12135 556 12201 559
rect 13383 556 13449 559
rect 14631 556 14697 559
rect 15879 556 15945 559
rect 17127 556 17193 559
rect 18375 556 18441 559
rect 19623 556 19689 559
rect 20871 556 20937 559
rect 22119 556 22185 559
rect 23367 556 23433 559
rect 24615 556 24681 559
rect 25863 556 25929 559
rect 27111 556 27177 559
rect 28359 556 28425 559
rect 29607 556 29673 559
rect 30855 556 30921 559
rect 32103 556 32169 559
rect 33351 556 33417 559
rect 34599 556 34665 559
rect 35847 556 35913 559
rect 37095 556 37161 559
rect 38343 556 38409 559
rect 39591 556 39657 559
rect 0 554 39936 556
rect 0 498 908 554
rect 964 498 2156 554
rect 2212 498 3404 554
rect 3460 498 4652 554
rect 4708 498 5900 554
rect 5956 498 7148 554
rect 7204 498 8396 554
rect 8452 498 9644 554
rect 9700 498 10892 554
rect 10948 498 12140 554
rect 12196 498 13388 554
rect 13444 498 14636 554
rect 14692 498 15884 554
rect 15940 498 17132 554
rect 17188 498 18380 554
rect 18436 498 19628 554
rect 19684 498 20876 554
rect 20932 498 22124 554
rect 22180 498 23372 554
rect 23428 498 24620 554
rect 24676 498 25868 554
rect 25924 498 27116 554
rect 27172 498 28364 554
rect 28420 498 29612 554
rect 29668 498 30860 554
rect 30916 498 32108 554
rect 32164 498 33356 554
rect 33412 498 34604 554
rect 34660 498 35852 554
rect 35908 498 37100 554
rect 37156 498 38348 554
rect 38404 498 39596 554
rect 39652 498 39936 554
rect 0 496 39936 498
rect 903 493 969 496
rect 2151 493 2217 496
rect 3399 493 3465 496
rect 4647 493 4713 496
rect 5895 493 5961 496
rect 7143 493 7209 496
rect 8391 493 8457 496
rect 9639 493 9705 496
rect 10887 493 10953 496
rect 12135 493 12201 496
rect 13383 493 13449 496
rect 14631 493 14697 496
rect 15879 493 15945 496
rect 17127 493 17193 496
rect 18375 493 18441 496
rect 19623 493 19689 496
rect 20871 493 20937 496
rect 22119 493 22185 496
rect 23367 493 23433 496
rect 24615 493 24681 496
rect 25863 493 25929 496
rect 27111 493 27177 496
rect 28359 493 28425 496
rect 29607 493 29673 496
rect 30855 493 30921 496
rect 32103 493 32169 496
rect 33351 493 33417 496
rect 34599 493 34665 496
rect 35847 493 35913 496
rect 37095 493 37161 496
rect 38343 493 38409 496
rect 39591 493 39657 496
rect 279 432 345 435
rect 1527 432 1593 435
rect 2775 432 2841 435
rect 4023 432 4089 435
rect 5271 432 5337 435
rect 6519 432 6585 435
rect 7767 432 7833 435
rect 9015 432 9081 435
rect 10263 432 10329 435
rect 11511 432 11577 435
rect 12759 432 12825 435
rect 14007 432 14073 435
rect 15255 432 15321 435
rect 16503 432 16569 435
rect 17751 432 17817 435
rect 18999 432 19065 435
rect 20247 432 20313 435
rect 21495 432 21561 435
rect 22743 432 22809 435
rect 23991 432 24057 435
rect 25239 432 25305 435
rect 26487 432 26553 435
rect 27735 432 27801 435
rect 28983 432 29049 435
rect 30231 432 30297 435
rect 31479 432 31545 435
rect 32727 432 32793 435
rect 33975 432 34041 435
rect 35223 432 35289 435
rect 36471 432 36537 435
rect 37719 432 37785 435
rect 38967 432 39033 435
rect 0 430 39936 432
rect 0 374 284 430
rect 340 374 1532 430
rect 1588 374 2780 430
rect 2836 374 4028 430
rect 4084 374 5276 430
rect 5332 374 6524 430
rect 6580 374 7772 430
rect 7828 374 9020 430
rect 9076 374 10268 430
rect 10324 374 11516 430
rect 11572 374 12764 430
rect 12820 374 14012 430
rect 14068 374 15260 430
rect 15316 374 16508 430
rect 16564 374 17756 430
rect 17812 374 19004 430
rect 19060 374 20252 430
rect 20308 374 21500 430
rect 21556 374 22748 430
rect 22804 374 23996 430
rect 24052 374 25244 430
rect 25300 374 26492 430
rect 26548 374 27740 430
rect 27796 374 28988 430
rect 29044 374 30236 430
rect 30292 374 31484 430
rect 31540 374 32732 430
rect 32788 374 33980 430
rect 34036 374 35228 430
rect 35284 374 36476 430
rect 36532 374 37724 430
rect 37780 374 38972 430
rect 39028 374 39936 430
rect 0 372 39936 374
rect 279 369 345 372
rect 1527 369 1593 372
rect 2775 369 2841 372
rect 4023 369 4089 372
rect 5271 369 5337 372
rect 6519 369 6585 372
rect 7767 369 7833 372
rect 9015 369 9081 372
rect 10263 369 10329 372
rect 11511 369 11577 372
rect 12759 369 12825 372
rect 14007 369 14073 372
rect 15255 369 15321 372
rect 16503 369 16569 372
rect 17751 369 17817 372
rect 18999 369 19065 372
rect 20247 369 20313 372
rect 21495 369 21561 372
rect 22743 369 22809 372
rect 23991 369 24057 372
rect 25239 369 25305 372
rect 26487 369 26553 372
rect 27735 369 27801 372
rect 28983 369 29049 372
rect 30231 369 30297 372
rect 31479 369 31545 372
rect 32727 369 32793 372
rect 33975 369 34041 372
rect 35223 369 35289 372
rect 36471 369 36537 372
rect 37719 369 37785 372
rect 38967 369 39033 372
rect 61 278 127 281
rect 1121 278 1187 281
rect 61 276 1187 278
rect 61 220 66 276
rect 122 220 1126 276
rect 1182 220 1187 276
rect 61 218 1187 220
rect 61 215 127 218
rect 1121 215 1187 218
rect 1309 278 1375 281
rect 2369 278 2435 281
rect 1309 276 2435 278
rect 1309 220 1314 276
rect 1370 220 2374 276
rect 2430 220 2435 276
rect 1309 218 2435 220
rect 1309 215 1375 218
rect 2369 215 2435 218
rect 2557 278 2623 281
rect 3617 278 3683 281
rect 2557 276 3683 278
rect 2557 220 2562 276
rect 2618 220 3622 276
rect 3678 220 3683 276
rect 2557 218 3683 220
rect 2557 215 2623 218
rect 3617 215 3683 218
rect 3805 278 3871 281
rect 4865 278 4931 281
rect 3805 276 4931 278
rect 3805 220 3810 276
rect 3866 220 4870 276
rect 4926 220 4931 276
rect 3805 218 4931 220
rect 3805 215 3871 218
rect 4865 215 4931 218
rect 5053 278 5119 281
rect 6113 278 6179 281
rect 5053 276 6179 278
rect 5053 220 5058 276
rect 5114 220 6118 276
rect 6174 220 6179 276
rect 5053 218 6179 220
rect 5053 215 5119 218
rect 6113 215 6179 218
rect 6301 278 6367 281
rect 7361 278 7427 281
rect 6301 276 7427 278
rect 6301 220 6306 276
rect 6362 220 7366 276
rect 7422 220 7427 276
rect 6301 218 7427 220
rect 6301 215 6367 218
rect 7361 215 7427 218
rect 7549 278 7615 281
rect 8609 278 8675 281
rect 7549 276 8675 278
rect 7549 220 7554 276
rect 7610 220 8614 276
rect 8670 220 8675 276
rect 7549 218 8675 220
rect 7549 215 7615 218
rect 8609 215 8675 218
rect 8797 278 8863 281
rect 9857 278 9923 281
rect 8797 276 9923 278
rect 8797 220 8802 276
rect 8858 220 9862 276
rect 9918 220 9923 276
rect 8797 218 9923 220
rect 8797 215 8863 218
rect 9857 215 9923 218
rect 10045 278 10111 281
rect 11105 278 11171 281
rect 10045 276 11171 278
rect 10045 220 10050 276
rect 10106 220 11110 276
rect 11166 220 11171 276
rect 10045 218 11171 220
rect 10045 215 10111 218
rect 11105 215 11171 218
rect 11293 278 11359 281
rect 12353 278 12419 281
rect 11293 276 12419 278
rect 11293 220 11298 276
rect 11354 220 12358 276
rect 12414 220 12419 276
rect 11293 218 12419 220
rect 11293 215 11359 218
rect 12353 215 12419 218
rect 12541 278 12607 281
rect 13601 278 13667 281
rect 12541 276 13667 278
rect 12541 220 12546 276
rect 12602 220 13606 276
rect 13662 220 13667 276
rect 12541 218 13667 220
rect 12541 215 12607 218
rect 13601 215 13667 218
rect 13789 278 13855 281
rect 14849 278 14915 281
rect 13789 276 14915 278
rect 13789 220 13794 276
rect 13850 220 14854 276
rect 14910 220 14915 276
rect 13789 218 14915 220
rect 13789 215 13855 218
rect 14849 215 14915 218
rect 15037 278 15103 281
rect 16097 278 16163 281
rect 15037 276 16163 278
rect 15037 220 15042 276
rect 15098 220 16102 276
rect 16158 220 16163 276
rect 15037 218 16163 220
rect 15037 215 15103 218
rect 16097 215 16163 218
rect 16285 278 16351 281
rect 17345 278 17411 281
rect 16285 276 17411 278
rect 16285 220 16290 276
rect 16346 220 17350 276
rect 17406 220 17411 276
rect 16285 218 17411 220
rect 16285 215 16351 218
rect 17345 215 17411 218
rect 17533 278 17599 281
rect 18593 278 18659 281
rect 17533 276 18659 278
rect 17533 220 17538 276
rect 17594 220 18598 276
rect 18654 220 18659 276
rect 17533 218 18659 220
rect 17533 215 17599 218
rect 18593 215 18659 218
rect 18781 278 18847 281
rect 19841 278 19907 281
rect 18781 276 19907 278
rect 18781 220 18786 276
rect 18842 220 19846 276
rect 19902 220 19907 276
rect 18781 218 19907 220
rect 18781 215 18847 218
rect 19841 215 19907 218
rect 20029 278 20095 281
rect 21089 278 21155 281
rect 20029 276 21155 278
rect 20029 220 20034 276
rect 20090 220 21094 276
rect 21150 220 21155 276
rect 20029 218 21155 220
rect 20029 215 20095 218
rect 21089 215 21155 218
rect 21277 278 21343 281
rect 22337 278 22403 281
rect 21277 276 22403 278
rect 21277 220 21282 276
rect 21338 220 22342 276
rect 22398 220 22403 276
rect 21277 218 22403 220
rect 21277 215 21343 218
rect 22337 215 22403 218
rect 22525 278 22591 281
rect 23585 278 23651 281
rect 22525 276 23651 278
rect 22525 220 22530 276
rect 22586 220 23590 276
rect 23646 220 23651 276
rect 22525 218 23651 220
rect 22525 215 22591 218
rect 23585 215 23651 218
rect 23773 278 23839 281
rect 24833 278 24899 281
rect 23773 276 24899 278
rect 23773 220 23778 276
rect 23834 220 24838 276
rect 24894 220 24899 276
rect 23773 218 24899 220
rect 23773 215 23839 218
rect 24833 215 24899 218
rect 25021 278 25087 281
rect 26081 278 26147 281
rect 25021 276 26147 278
rect 25021 220 25026 276
rect 25082 220 26086 276
rect 26142 220 26147 276
rect 25021 218 26147 220
rect 25021 215 25087 218
rect 26081 215 26147 218
rect 26269 278 26335 281
rect 27329 278 27395 281
rect 26269 276 27395 278
rect 26269 220 26274 276
rect 26330 220 27334 276
rect 27390 220 27395 276
rect 26269 218 27395 220
rect 26269 215 26335 218
rect 27329 215 27395 218
rect 27517 278 27583 281
rect 28577 278 28643 281
rect 27517 276 28643 278
rect 27517 220 27522 276
rect 27578 220 28582 276
rect 28638 220 28643 276
rect 27517 218 28643 220
rect 27517 215 27583 218
rect 28577 215 28643 218
rect 28765 278 28831 281
rect 29825 278 29891 281
rect 28765 276 29891 278
rect 28765 220 28770 276
rect 28826 220 29830 276
rect 29886 220 29891 276
rect 28765 218 29891 220
rect 28765 215 28831 218
rect 29825 215 29891 218
rect 30013 278 30079 281
rect 31073 278 31139 281
rect 30013 276 31139 278
rect 30013 220 30018 276
rect 30074 220 31078 276
rect 31134 220 31139 276
rect 30013 218 31139 220
rect 30013 215 30079 218
rect 31073 215 31139 218
rect 31261 278 31327 281
rect 32321 278 32387 281
rect 31261 276 32387 278
rect 31261 220 31266 276
rect 31322 220 32326 276
rect 32382 220 32387 276
rect 31261 218 32387 220
rect 31261 215 31327 218
rect 32321 215 32387 218
rect 32509 278 32575 281
rect 33569 278 33635 281
rect 32509 276 33635 278
rect 32509 220 32514 276
rect 32570 220 33574 276
rect 33630 220 33635 276
rect 32509 218 33635 220
rect 32509 215 32575 218
rect 33569 215 33635 218
rect 33757 278 33823 281
rect 34817 278 34883 281
rect 33757 276 34883 278
rect 33757 220 33762 276
rect 33818 220 34822 276
rect 34878 220 34883 276
rect 33757 218 34883 220
rect 33757 215 33823 218
rect 34817 215 34883 218
rect 35005 278 35071 281
rect 36065 278 36131 281
rect 35005 276 36131 278
rect 35005 220 35010 276
rect 35066 220 36070 276
rect 36126 220 36131 276
rect 35005 218 36131 220
rect 35005 215 35071 218
rect 36065 215 36131 218
rect 36253 278 36319 281
rect 37313 278 37379 281
rect 36253 276 37379 278
rect 36253 220 36258 276
rect 36314 220 37318 276
rect 37374 220 37379 276
rect 36253 218 37379 220
rect 36253 215 36319 218
rect 37313 215 37379 218
rect 37501 278 37567 281
rect 38561 278 38627 281
rect 37501 276 38627 278
rect 37501 220 37506 276
rect 37562 220 38566 276
rect 38622 220 38627 276
rect 37501 218 38627 220
rect 37501 215 37567 218
rect 38561 215 38627 218
rect 38749 278 38815 281
rect 39809 278 39875 281
rect 38749 276 39875 278
rect 38749 220 38754 276
rect 38810 220 39814 276
rect 39870 220 39875 276
rect 38749 218 39875 220
rect 38749 215 38815 218
rect 39809 215 39875 218
rect 525 154 591 157
rect 657 154 723 157
rect 525 152 723 154
rect 525 96 530 152
rect 586 96 662 152
rect 718 96 723 152
rect 525 94 723 96
rect 525 91 591 94
rect 657 91 723 94
rect 1773 154 1839 157
rect 1905 154 1971 157
rect 1773 152 1971 154
rect 1773 96 1778 152
rect 1834 96 1910 152
rect 1966 96 1971 152
rect 1773 94 1971 96
rect 1773 91 1839 94
rect 1905 91 1971 94
rect 3021 154 3087 157
rect 3153 154 3219 157
rect 3021 152 3219 154
rect 3021 96 3026 152
rect 3082 96 3158 152
rect 3214 96 3219 152
rect 3021 94 3219 96
rect 3021 91 3087 94
rect 3153 91 3219 94
rect 4269 154 4335 157
rect 4401 154 4467 157
rect 4269 152 4467 154
rect 4269 96 4274 152
rect 4330 96 4406 152
rect 4462 96 4467 152
rect 4269 94 4467 96
rect 4269 91 4335 94
rect 4401 91 4467 94
rect 5517 154 5583 157
rect 5649 154 5715 157
rect 5517 152 5715 154
rect 5517 96 5522 152
rect 5578 96 5654 152
rect 5710 96 5715 152
rect 5517 94 5715 96
rect 5517 91 5583 94
rect 5649 91 5715 94
rect 6765 154 6831 157
rect 6897 154 6963 157
rect 6765 152 6963 154
rect 6765 96 6770 152
rect 6826 96 6902 152
rect 6958 96 6963 152
rect 6765 94 6963 96
rect 6765 91 6831 94
rect 6897 91 6963 94
rect 8013 154 8079 157
rect 8145 154 8211 157
rect 8013 152 8211 154
rect 8013 96 8018 152
rect 8074 96 8150 152
rect 8206 96 8211 152
rect 8013 94 8211 96
rect 8013 91 8079 94
rect 8145 91 8211 94
rect 9261 154 9327 157
rect 9393 154 9459 157
rect 9261 152 9459 154
rect 9261 96 9266 152
rect 9322 96 9398 152
rect 9454 96 9459 152
rect 9261 94 9459 96
rect 9261 91 9327 94
rect 9393 91 9459 94
rect 10509 154 10575 157
rect 10641 154 10707 157
rect 10509 152 10707 154
rect 10509 96 10514 152
rect 10570 96 10646 152
rect 10702 96 10707 152
rect 10509 94 10707 96
rect 10509 91 10575 94
rect 10641 91 10707 94
rect 11757 154 11823 157
rect 11889 154 11955 157
rect 11757 152 11955 154
rect 11757 96 11762 152
rect 11818 96 11894 152
rect 11950 96 11955 152
rect 11757 94 11955 96
rect 11757 91 11823 94
rect 11889 91 11955 94
rect 13005 154 13071 157
rect 13137 154 13203 157
rect 13005 152 13203 154
rect 13005 96 13010 152
rect 13066 96 13142 152
rect 13198 96 13203 152
rect 13005 94 13203 96
rect 13005 91 13071 94
rect 13137 91 13203 94
rect 14253 154 14319 157
rect 14385 154 14451 157
rect 14253 152 14451 154
rect 14253 96 14258 152
rect 14314 96 14390 152
rect 14446 96 14451 152
rect 14253 94 14451 96
rect 14253 91 14319 94
rect 14385 91 14451 94
rect 15501 154 15567 157
rect 15633 154 15699 157
rect 15501 152 15699 154
rect 15501 96 15506 152
rect 15562 96 15638 152
rect 15694 96 15699 152
rect 15501 94 15699 96
rect 15501 91 15567 94
rect 15633 91 15699 94
rect 16749 154 16815 157
rect 16881 154 16947 157
rect 16749 152 16947 154
rect 16749 96 16754 152
rect 16810 96 16886 152
rect 16942 96 16947 152
rect 16749 94 16947 96
rect 16749 91 16815 94
rect 16881 91 16947 94
rect 17997 154 18063 157
rect 18129 154 18195 157
rect 17997 152 18195 154
rect 17997 96 18002 152
rect 18058 96 18134 152
rect 18190 96 18195 152
rect 17997 94 18195 96
rect 17997 91 18063 94
rect 18129 91 18195 94
rect 19245 154 19311 157
rect 19377 154 19443 157
rect 19245 152 19443 154
rect 19245 96 19250 152
rect 19306 96 19382 152
rect 19438 96 19443 152
rect 19245 94 19443 96
rect 19245 91 19311 94
rect 19377 91 19443 94
rect 20493 154 20559 157
rect 20625 154 20691 157
rect 20493 152 20691 154
rect 20493 96 20498 152
rect 20554 96 20630 152
rect 20686 96 20691 152
rect 20493 94 20691 96
rect 20493 91 20559 94
rect 20625 91 20691 94
rect 21741 154 21807 157
rect 21873 154 21939 157
rect 21741 152 21939 154
rect 21741 96 21746 152
rect 21802 96 21878 152
rect 21934 96 21939 152
rect 21741 94 21939 96
rect 21741 91 21807 94
rect 21873 91 21939 94
rect 22989 154 23055 157
rect 23121 154 23187 157
rect 22989 152 23187 154
rect 22989 96 22994 152
rect 23050 96 23126 152
rect 23182 96 23187 152
rect 22989 94 23187 96
rect 22989 91 23055 94
rect 23121 91 23187 94
rect 24237 154 24303 157
rect 24369 154 24435 157
rect 24237 152 24435 154
rect 24237 96 24242 152
rect 24298 96 24374 152
rect 24430 96 24435 152
rect 24237 94 24435 96
rect 24237 91 24303 94
rect 24369 91 24435 94
rect 25485 154 25551 157
rect 25617 154 25683 157
rect 25485 152 25683 154
rect 25485 96 25490 152
rect 25546 96 25622 152
rect 25678 96 25683 152
rect 25485 94 25683 96
rect 25485 91 25551 94
rect 25617 91 25683 94
rect 26733 154 26799 157
rect 26865 154 26931 157
rect 26733 152 26931 154
rect 26733 96 26738 152
rect 26794 96 26870 152
rect 26926 96 26931 152
rect 26733 94 26931 96
rect 26733 91 26799 94
rect 26865 91 26931 94
rect 27981 154 28047 157
rect 28113 154 28179 157
rect 27981 152 28179 154
rect 27981 96 27986 152
rect 28042 96 28118 152
rect 28174 96 28179 152
rect 27981 94 28179 96
rect 27981 91 28047 94
rect 28113 91 28179 94
rect 29229 154 29295 157
rect 29361 154 29427 157
rect 29229 152 29427 154
rect 29229 96 29234 152
rect 29290 96 29366 152
rect 29422 96 29427 152
rect 29229 94 29427 96
rect 29229 91 29295 94
rect 29361 91 29427 94
rect 30477 154 30543 157
rect 30609 154 30675 157
rect 30477 152 30675 154
rect 30477 96 30482 152
rect 30538 96 30614 152
rect 30670 96 30675 152
rect 30477 94 30675 96
rect 30477 91 30543 94
rect 30609 91 30675 94
rect 31725 154 31791 157
rect 31857 154 31923 157
rect 31725 152 31923 154
rect 31725 96 31730 152
rect 31786 96 31862 152
rect 31918 96 31923 152
rect 31725 94 31923 96
rect 31725 91 31791 94
rect 31857 91 31923 94
rect 32973 154 33039 157
rect 33105 154 33171 157
rect 32973 152 33171 154
rect 32973 96 32978 152
rect 33034 96 33110 152
rect 33166 96 33171 152
rect 32973 94 33171 96
rect 32973 91 33039 94
rect 33105 91 33171 94
rect 34221 154 34287 157
rect 34353 154 34419 157
rect 34221 152 34419 154
rect 34221 96 34226 152
rect 34282 96 34358 152
rect 34414 96 34419 152
rect 34221 94 34419 96
rect 34221 91 34287 94
rect 34353 91 34419 94
rect 35469 154 35535 157
rect 35601 154 35667 157
rect 35469 152 35667 154
rect 35469 96 35474 152
rect 35530 96 35606 152
rect 35662 96 35667 152
rect 35469 94 35667 96
rect 35469 91 35535 94
rect 35601 91 35667 94
rect 36717 154 36783 157
rect 36849 154 36915 157
rect 36717 152 36915 154
rect 36717 96 36722 152
rect 36778 96 36854 152
rect 36910 96 36915 152
rect 36717 94 36915 96
rect 36717 91 36783 94
rect 36849 91 36915 94
rect 37965 154 38031 157
rect 38097 154 38163 157
rect 37965 152 38163 154
rect 37965 96 37970 152
rect 38026 96 38102 152
rect 38158 96 38163 152
rect 37965 94 38163 96
rect 37965 91 38031 94
rect 38097 91 38163 94
rect 39213 154 39279 157
rect 39345 154 39411 157
rect 39213 152 39411 154
rect 39213 96 39218 152
rect 39274 96 39350 152
rect 39406 96 39411 152
rect 39213 94 39411 96
rect 39213 91 39279 94
rect 39345 91 39411 94
use contact_19  contact_19_0
timestamp 1683767628
transform 1 0 4023 0 1 369
box 0 0 1 1
use contact_19  contact_19_1
timestamp 1683767628
transform 1 0 279 0 1 369
box 0 0 1 1
use contact_19  contact_19_2
timestamp 1683767628
transform 1 0 2775 0 1 369
box 0 0 1 1
use contact_19  contact_19_3
timestamp 1683767628
transform 1 0 1527 0 1 369
box 0 0 1 1
use contact_19  contact_19_4
timestamp 1683767628
transform 1 0 4647 0 1 493
box 0 0 1 1
use contact_19  contact_19_5
timestamp 1683767628
transform 1 0 3399 0 1 493
box 0 0 1 1
use contact_19  contact_19_6
timestamp 1683767628
transform 1 0 2151 0 1 493
box 0 0 1 1
use contact_19  contact_19_7
timestamp 1683767628
transform 1 0 903 0 1 493
box 0 0 1 1
use contact_19  contact_19_8
timestamp 1683767628
transform 1 0 9015 0 1 369
box 0 0 1 1
use contact_19  contact_19_9
timestamp 1683767628
transform 1 0 7767 0 1 369
box 0 0 1 1
use contact_19  contact_19_10
timestamp 1683767628
transform 1 0 6519 0 1 369
box 0 0 1 1
use contact_19  contact_19_11
timestamp 1683767628
transform 1 0 5271 0 1 369
box 0 0 1 1
use contact_19  contact_19_12
timestamp 1683767628
transform 1 0 9639 0 1 493
box 0 0 1 1
use contact_19  contact_19_13
timestamp 1683767628
transform 1 0 8391 0 1 493
box 0 0 1 1
use contact_19  contact_19_14
timestamp 1683767628
transform 1 0 7143 0 1 493
box 0 0 1 1
use contact_19  contact_19_15
timestamp 1683767628
transform 1 0 5895 0 1 493
box 0 0 1 1
use contact_19  contact_19_16
timestamp 1683767628
transform 1 0 14007 0 1 369
box 0 0 1 1
use contact_19  contact_19_17
timestamp 1683767628
transform 1 0 10263 0 1 369
box 0 0 1 1
use contact_19  contact_19_18
timestamp 1683767628
transform 1 0 12759 0 1 369
box 0 0 1 1
use contact_19  contact_19_19
timestamp 1683767628
transform 1 0 11511 0 1 369
box 0 0 1 1
use contact_19  contact_19_20
timestamp 1683767628
transform 1 0 14631 0 1 493
box 0 0 1 1
use contact_19  contact_19_21
timestamp 1683767628
transform 1 0 13383 0 1 493
box 0 0 1 1
use contact_19  contact_19_22
timestamp 1683767628
transform 1 0 12135 0 1 493
box 0 0 1 1
use contact_19  contact_19_23
timestamp 1683767628
transform 1 0 10887 0 1 493
box 0 0 1 1
use contact_19  contact_19_24
timestamp 1683767628
transform 1 0 18999 0 1 369
box 0 0 1 1
use contact_19  contact_19_25
timestamp 1683767628
transform 1 0 17751 0 1 369
box 0 0 1 1
use contact_19  contact_19_26
timestamp 1683767628
transform 1 0 16503 0 1 369
box 0 0 1 1
use contact_19  contact_19_27
timestamp 1683767628
transform 1 0 15255 0 1 369
box 0 0 1 1
use contact_19  contact_19_28
timestamp 1683767628
transform 1 0 19623 0 1 493
box 0 0 1 1
use contact_19  contact_19_29
timestamp 1683767628
transform 1 0 18375 0 1 493
box 0 0 1 1
use contact_19  contact_19_30
timestamp 1683767628
transform 1 0 17127 0 1 493
box 0 0 1 1
use contact_19  contact_19_31
timestamp 1683767628
transform 1 0 15879 0 1 493
box 0 0 1 1
use contact_19  contact_19_32
timestamp 1683767628
transform 1 0 23991 0 1 369
box 0 0 1 1
use contact_19  contact_19_33
timestamp 1683767628
transform 1 0 20247 0 1 369
box 0 0 1 1
use contact_19  contact_19_34
timestamp 1683767628
transform 1 0 22743 0 1 369
box 0 0 1 1
use contact_19  contact_19_35
timestamp 1683767628
transform 1 0 21495 0 1 369
box 0 0 1 1
use contact_19  contact_19_36
timestamp 1683767628
transform 1 0 24615 0 1 493
box 0 0 1 1
use contact_19  contact_19_37
timestamp 1683767628
transform 1 0 23367 0 1 493
box 0 0 1 1
use contact_19  contact_19_38
timestamp 1683767628
transform 1 0 22119 0 1 493
box 0 0 1 1
use contact_19  contact_19_39
timestamp 1683767628
transform 1 0 20871 0 1 493
box 0 0 1 1
use contact_19  contact_19_40
timestamp 1683767628
transform 1 0 28983 0 1 369
box 0 0 1 1
use contact_19  contact_19_41
timestamp 1683767628
transform 1 0 27735 0 1 369
box 0 0 1 1
use contact_19  contact_19_42
timestamp 1683767628
transform 1 0 26487 0 1 369
box 0 0 1 1
use contact_19  contact_19_43
timestamp 1683767628
transform 1 0 25239 0 1 369
box 0 0 1 1
use contact_19  contact_19_44
timestamp 1683767628
transform 1 0 29607 0 1 493
box 0 0 1 1
use contact_19  contact_19_45
timestamp 1683767628
transform 1 0 28359 0 1 493
box 0 0 1 1
use contact_19  contact_19_46
timestamp 1683767628
transform 1 0 27111 0 1 493
box 0 0 1 1
use contact_19  contact_19_47
timestamp 1683767628
transform 1 0 25863 0 1 493
box 0 0 1 1
use contact_19  contact_19_48
timestamp 1683767628
transform 1 0 30231 0 1 369
box 0 0 1 1
use contact_19  contact_19_49
timestamp 1683767628
transform 1 0 32727 0 1 369
box 0 0 1 1
use contact_19  contact_19_50
timestamp 1683767628
transform 1 0 31479 0 1 369
box 0 0 1 1
use contact_19  contact_19_51
timestamp 1683767628
transform 1 0 34599 0 1 493
box 0 0 1 1
use contact_19  contact_19_52
timestamp 1683767628
transform 1 0 33351 0 1 493
box 0 0 1 1
use contact_19  contact_19_53
timestamp 1683767628
transform 1 0 32103 0 1 493
box 0 0 1 1
use contact_19  contact_19_54
timestamp 1683767628
transform 1 0 30855 0 1 493
box 0 0 1 1
use contact_19  contact_19_55
timestamp 1683767628
transform 1 0 33975 0 1 369
box 0 0 1 1
use contact_19  contact_19_56
timestamp 1683767628
transform 1 0 38967 0 1 369
box 0 0 1 1
use contact_19  contact_19_57
timestamp 1683767628
transform 1 0 37719 0 1 369
box 0 0 1 1
use contact_19  contact_19_58
timestamp 1683767628
transform 1 0 36471 0 1 369
box 0 0 1 1
use contact_19  contact_19_59
timestamp 1683767628
transform 1 0 35223 0 1 369
box 0 0 1 1
use contact_19  contact_19_60
timestamp 1683767628
transform 1 0 39591 0 1 493
box 0 0 1 1
use contact_19  contact_19_61
timestamp 1683767628
transform 1 0 38343 0 1 493
box 0 0 1 1
use contact_19  contact_19_62
timestamp 1683767628
transform 1 0 37095 0 1 493
box 0 0 1 1
use contact_19  contact_19_63
timestamp 1683767628
transform 1 0 35847 0 1 493
box 0 0 1 1
use contact_20  contact_20_0
timestamp 1683767628
transform 1 0 283 0 1 369
box 0 0 1 1
use contact_20  contact_20_1
timestamp 1683767628
transform 1 0 4651 0 1 493
box 0 0 1 1
use contact_20  contact_20_2
timestamp 1683767628
transform 1 0 4027 0 1 369
box 0 0 1 1
use contact_20  contact_20_3
timestamp 1683767628
transform 1 0 907 0 1 493
box 0 0 1 1
use contact_20  contact_20_4
timestamp 1683767628
transform 1 0 3403 0 1 493
box 0 0 1 1
use contact_20  contact_20_5
timestamp 1683767628
transform 1 0 2779 0 1 369
box 0 0 1 1
use contact_20  contact_20_6
timestamp 1683767628
transform 1 0 2155 0 1 493
box 0 0 1 1
use contact_20  contact_20_7
timestamp 1683767628
transform 1 0 1531 0 1 369
box 0 0 1 1
use contact_20  contact_20_8
timestamp 1683767628
transform 1 0 9643 0 1 493
box 0 0 1 1
use contact_20  contact_20_9
timestamp 1683767628
transform 1 0 9019 0 1 369
box 0 0 1 1
use contact_20  contact_20_10
timestamp 1683767628
transform 1 0 8395 0 1 493
box 0 0 1 1
use contact_20  contact_20_11
timestamp 1683767628
transform 1 0 7771 0 1 369
box 0 0 1 1
use contact_20  contact_20_12
timestamp 1683767628
transform 1 0 7147 0 1 493
box 0 0 1 1
use contact_20  contact_20_13
timestamp 1683767628
transform 1 0 6523 0 1 369
box 0 0 1 1
use contact_20  contact_20_14
timestamp 1683767628
transform 1 0 5899 0 1 493
box 0 0 1 1
use contact_20  contact_20_15
timestamp 1683767628
transform 1 0 5275 0 1 369
box 0 0 1 1
use contact_20  contact_20_16
timestamp 1683767628
transform 1 0 10267 0 1 369
box 0 0 1 1
use contact_20  contact_20_17
timestamp 1683767628
transform 1 0 14635 0 1 493
box 0 0 1 1
use contact_20  contact_20_18
timestamp 1683767628
transform 1 0 14011 0 1 369
box 0 0 1 1
use contact_20  contact_20_19
timestamp 1683767628
transform 1 0 10891 0 1 493
box 0 0 1 1
use contact_20  contact_20_20
timestamp 1683767628
transform 1 0 13387 0 1 493
box 0 0 1 1
use contact_20  contact_20_21
timestamp 1683767628
transform 1 0 12763 0 1 369
box 0 0 1 1
use contact_20  contact_20_22
timestamp 1683767628
transform 1 0 12139 0 1 493
box 0 0 1 1
use contact_20  contact_20_23
timestamp 1683767628
transform 1 0 11515 0 1 369
box 0 0 1 1
use contact_20  contact_20_24
timestamp 1683767628
transform 1 0 19627 0 1 493
box 0 0 1 1
use contact_20  contact_20_25
timestamp 1683767628
transform 1 0 19003 0 1 369
box 0 0 1 1
use contact_20  contact_20_26
timestamp 1683767628
transform 1 0 18379 0 1 493
box 0 0 1 1
use contact_20  contact_20_27
timestamp 1683767628
transform 1 0 17755 0 1 369
box 0 0 1 1
use contact_20  contact_20_28
timestamp 1683767628
transform 1 0 17131 0 1 493
box 0 0 1 1
use contact_20  contact_20_29
timestamp 1683767628
transform 1 0 16507 0 1 369
box 0 0 1 1
use contact_20  contact_20_30
timestamp 1683767628
transform 1 0 15883 0 1 493
box 0 0 1 1
use contact_20  contact_20_31
timestamp 1683767628
transform 1 0 15259 0 1 369
box 0 0 1 1
use contact_20  contact_20_32
timestamp 1683767628
transform 1 0 20251 0 1 369
box 0 0 1 1
use contact_20  contact_20_33
timestamp 1683767628
transform 1 0 24619 0 1 493
box 0 0 1 1
use contact_20  contact_20_34
timestamp 1683767628
transform 1 0 23995 0 1 369
box 0 0 1 1
use contact_20  contact_20_35
timestamp 1683767628
transform 1 0 20875 0 1 493
box 0 0 1 1
use contact_20  contact_20_36
timestamp 1683767628
transform 1 0 23371 0 1 493
box 0 0 1 1
use contact_20  contact_20_37
timestamp 1683767628
transform 1 0 22747 0 1 369
box 0 0 1 1
use contact_20  contact_20_38
timestamp 1683767628
transform 1 0 22123 0 1 493
box 0 0 1 1
use contact_20  contact_20_39
timestamp 1683767628
transform 1 0 21499 0 1 369
box 0 0 1 1
use contact_20  contact_20_40
timestamp 1683767628
transform 1 0 29611 0 1 493
box 0 0 1 1
use contact_20  contact_20_41
timestamp 1683767628
transform 1 0 28987 0 1 369
box 0 0 1 1
use contact_20  contact_20_42
timestamp 1683767628
transform 1 0 28363 0 1 493
box 0 0 1 1
use contact_20  contact_20_43
timestamp 1683767628
transform 1 0 27739 0 1 369
box 0 0 1 1
use contact_20  contact_20_44
timestamp 1683767628
transform 1 0 27115 0 1 493
box 0 0 1 1
use contact_20  contact_20_45
timestamp 1683767628
transform 1 0 26491 0 1 369
box 0 0 1 1
use contact_20  contact_20_46
timestamp 1683767628
transform 1 0 25867 0 1 493
box 0 0 1 1
use contact_20  contact_20_47
timestamp 1683767628
transform 1 0 25243 0 1 369
box 0 0 1 1
use contact_20  contact_20_48
timestamp 1683767628
transform 1 0 30859 0 1 493
box 0 0 1 1
use contact_20  contact_20_49
timestamp 1683767628
transform 1 0 33355 0 1 493
box 0 0 1 1
use contact_20  contact_20_50
timestamp 1683767628
transform 1 0 32731 0 1 369
box 0 0 1 1
use contact_20  contact_20_51
timestamp 1683767628
transform 1 0 32107 0 1 493
box 0 0 1 1
use contact_20  contact_20_52
timestamp 1683767628
transform 1 0 31483 0 1 369
box 0 0 1 1
use contact_20  contact_20_53
timestamp 1683767628
transform 1 0 30235 0 1 369
box 0 0 1 1
use contact_20  contact_20_54
timestamp 1683767628
transform 1 0 34603 0 1 493
box 0 0 1 1
use contact_20  contact_20_55
timestamp 1683767628
transform 1 0 33979 0 1 369
box 0 0 1 1
use contact_20  contact_20_56
timestamp 1683767628
transform 1 0 39595 0 1 493
box 0 0 1 1
use contact_20  contact_20_57
timestamp 1683767628
transform 1 0 38971 0 1 369
box 0 0 1 1
use contact_20  contact_20_58
timestamp 1683767628
transform 1 0 38347 0 1 493
box 0 0 1 1
use contact_20  contact_20_59
timestamp 1683767628
transform 1 0 37723 0 1 369
box 0 0 1 1
use contact_20  contact_20_60
timestamp 1683767628
transform 1 0 37099 0 1 493
box 0 0 1 1
use contact_20  contact_20_61
timestamp 1683767628
transform 1 0 36475 0 1 369
box 0 0 1 1
use contact_20  contact_20_62
timestamp 1683767628
transform 1 0 35851 0 1 493
box 0 0 1 1
use contact_20  contact_20_63
timestamp 1683767628
transform 1 0 35227 0 1 369
box 0 0 1 1
use contact_21  contact_21_0
timestamp 1683767628
transform 1 0 4648 0 1 494
box 0 0 1 1
use contact_21  contact_21_1
timestamp 1683767628
transform 1 0 904 0 1 494
box 0 0 1 1
use contact_21  contact_21_2
timestamp 1683767628
transform 1 0 4024 0 1 370
box 0 0 1 1
use contact_21  contact_21_3
timestamp 1683767628
transform 1 0 3400 0 1 494
box 0 0 1 1
use contact_21  contact_21_4
timestamp 1683767628
transform 1 0 2776 0 1 370
box 0 0 1 1
use contact_21  contact_21_5
timestamp 1683767628
transform 1 0 2152 0 1 494
box 0 0 1 1
use contact_21  contact_21_6
timestamp 1683767628
transform 1 0 1528 0 1 370
box 0 0 1 1
use contact_21  contact_21_7
timestamp 1683767628
transform 1 0 280 0 1 370
box 0 0 1 1
use contact_21  contact_21_8
timestamp 1683767628
transform 1 0 4402 0 1 92
box 0 0 1 1
use contact_21  contact_21_9
timestamp 1683767628
transform 1 0 4866 0 1 216
box 0 0 1 1
use contact_21  contact_21_10
timestamp 1683767628
transform 1 0 4270 0 1 92
box 0 0 1 1
use contact_21  contact_21_11
timestamp 1683767628
transform 1 0 3806 0 1 216
box 0 0 1 1
use contact_21  contact_21_12
timestamp 1683767628
transform 1 0 3154 0 1 92
box 0 0 1 1
use contact_21  contact_21_13
timestamp 1683767628
transform 1 0 3618 0 1 216
box 0 0 1 1
use contact_21  contact_21_14
timestamp 1683767628
transform 1 0 3022 0 1 92
box 0 0 1 1
use contact_21  contact_21_15
timestamp 1683767628
transform 1 0 2558 0 1 216
box 0 0 1 1
use contact_21  contact_21_16
timestamp 1683767628
transform 1 0 1906 0 1 92
box 0 0 1 1
use contact_21  contact_21_17
timestamp 1683767628
transform 1 0 2370 0 1 216
box 0 0 1 1
use contact_21  contact_21_18
timestamp 1683767628
transform 1 0 1774 0 1 92
box 0 0 1 1
use contact_21  contact_21_19
timestamp 1683767628
transform 1 0 1310 0 1 216
box 0 0 1 1
use contact_21  contact_21_20
timestamp 1683767628
transform 1 0 658 0 1 92
box 0 0 1 1
use contact_21  contact_21_21
timestamp 1683767628
transform 1 0 1122 0 1 216
box 0 0 1 1
use contact_21  contact_21_22
timestamp 1683767628
transform 1 0 526 0 1 92
box 0 0 1 1
use contact_21  contact_21_23
timestamp 1683767628
transform 1 0 62 0 1 216
box 0 0 1 1
use contact_21  contact_21_24
timestamp 1683767628
transform 1 0 9640 0 1 494
box 0 0 1 1
use contact_21  contact_21_25
timestamp 1683767628
transform 1 0 9016 0 1 370
box 0 0 1 1
use contact_21  contact_21_26
timestamp 1683767628
transform 1 0 8392 0 1 494
box 0 0 1 1
use contact_21  contact_21_27
timestamp 1683767628
transform 1 0 7768 0 1 370
box 0 0 1 1
use contact_21  contact_21_28
timestamp 1683767628
transform 1 0 7144 0 1 494
box 0 0 1 1
use contact_21  contact_21_29
timestamp 1683767628
transform 1 0 6520 0 1 370
box 0 0 1 1
use contact_21  contact_21_30
timestamp 1683767628
transform 1 0 5896 0 1 494
box 0 0 1 1
use contact_21  contact_21_31
timestamp 1683767628
transform 1 0 5272 0 1 370
box 0 0 1 1
use contact_21  contact_21_32
timestamp 1683767628
transform 1 0 9394 0 1 92
box 0 0 1 1
use contact_21  contact_21_33
timestamp 1683767628
transform 1 0 9858 0 1 216
box 0 0 1 1
use contact_21  contact_21_34
timestamp 1683767628
transform 1 0 9262 0 1 92
box 0 0 1 1
use contact_21  contact_21_35
timestamp 1683767628
transform 1 0 8798 0 1 216
box 0 0 1 1
use contact_21  contact_21_36
timestamp 1683767628
transform 1 0 8146 0 1 92
box 0 0 1 1
use contact_21  contact_21_37
timestamp 1683767628
transform 1 0 8610 0 1 216
box 0 0 1 1
use contact_21  contact_21_38
timestamp 1683767628
transform 1 0 8014 0 1 92
box 0 0 1 1
use contact_21  contact_21_39
timestamp 1683767628
transform 1 0 7550 0 1 216
box 0 0 1 1
use contact_21  contact_21_40
timestamp 1683767628
transform 1 0 6898 0 1 92
box 0 0 1 1
use contact_21  contact_21_41
timestamp 1683767628
transform 1 0 7362 0 1 216
box 0 0 1 1
use contact_21  contact_21_42
timestamp 1683767628
transform 1 0 6766 0 1 92
box 0 0 1 1
use contact_21  contact_21_43
timestamp 1683767628
transform 1 0 6302 0 1 216
box 0 0 1 1
use contact_21  contact_21_44
timestamp 1683767628
transform 1 0 5650 0 1 92
box 0 0 1 1
use contact_21  contact_21_45
timestamp 1683767628
transform 1 0 6114 0 1 216
box 0 0 1 1
use contact_21  contact_21_46
timestamp 1683767628
transform 1 0 5518 0 1 92
box 0 0 1 1
use contact_21  contact_21_47
timestamp 1683767628
transform 1 0 5054 0 1 216
box 0 0 1 1
use contact_21  contact_21_48
timestamp 1683767628
transform 1 0 14386 0 1 92
box 0 0 1 1
use contact_21  contact_21_49
timestamp 1683767628
transform 1 0 14850 0 1 216
box 0 0 1 1
use contact_21  contact_21_50
timestamp 1683767628
transform 1 0 14254 0 1 92
box 0 0 1 1
use contact_21  contact_21_51
timestamp 1683767628
transform 1 0 13790 0 1 216
box 0 0 1 1
use contact_21  contact_21_52
timestamp 1683767628
transform 1 0 13138 0 1 92
box 0 0 1 1
use contact_21  contact_21_53
timestamp 1683767628
transform 1 0 13602 0 1 216
box 0 0 1 1
use contact_21  contact_21_54
timestamp 1683767628
transform 1 0 13006 0 1 92
box 0 0 1 1
use contact_21  contact_21_55
timestamp 1683767628
transform 1 0 12542 0 1 216
box 0 0 1 1
use contact_21  contact_21_56
timestamp 1683767628
transform 1 0 11890 0 1 92
box 0 0 1 1
use contact_21  contact_21_57
timestamp 1683767628
transform 1 0 12354 0 1 216
box 0 0 1 1
use contact_21  contact_21_58
timestamp 1683767628
transform 1 0 11758 0 1 92
box 0 0 1 1
use contact_21  contact_21_59
timestamp 1683767628
transform 1 0 11294 0 1 216
box 0 0 1 1
use contact_21  contact_21_60
timestamp 1683767628
transform 1 0 10642 0 1 92
box 0 0 1 1
use contact_21  contact_21_61
timestamp 1683767628
transform 1 0 11106 0 1 216
box 0 0 1 1
use contact_21  contact_21_62
timestamp 1683767628
transform 1 0 10510 0 1 92
box 0 0 1 1
use contact_21  contact_21_63
timestamp 1683767628
transform 1 0 10046 0 1 216
box 0 0 1 1
use contact_21  contact_21_64
timestamp 1683767628
transform 1 0 14632 0 1 494
box 0 0 1 1
use contact_21  contact_21_65
timestamp 1683767628
transform 1 0 10888 0 1 494
box 0 0 1 1
use contact_21  contact_21_66
timestamp 1683767628
transform 1 0 14008 0 1 370
box 0 0 1 1
use contact_21  contact_21_67
timestamp 1683767628
transform 1 0 13384 0 1 494
box 0 0 1 1
use contact_21  contact_21_68
timestamp 1683767628
transform 1 0 12760 0 1 370
box 0 0 1 1
use contact_21  contact_21_69
timestamp 1683767628
transform 1 0 12136 0 1 494
box 0 0 1 1
use contact_21  contact_21_70
timestamp 1683767628
transform 1 0 11512 0 1 370
box 0 0 1 1
use contact_21  contact_21_71
timestamp 1683767628
transform 1 0 10264 0 1 370
box 0 0 1 1
use contact_21  contact_21_72
timestamp 1683767628
transform 1 0 19624 0 1 494
box 0 0 1 1
use contact_21  contact_21_73
timestamp 1683767628
transform 1 0 19000 0 1 370
box 0 0 1 1
use contact_21  contact_21_74
timestamp 1683767628
transform 1 0 18376 0 1 494
box 0 0 1 1
use contact_21  contact_21_75
timestamp 1683767628
transform 1 0 17752 0 1 370
box 0 0 1 1
use contact_21  contact_21_76
timestamp 1683767628
transform 1 0 17128 0 1 494
box 0 0 1 1
use contact_21  contact_21_77
timestamp 1683767628
transform 1 0 16504 0 1 370
box 0 0 1 1
use contact_21  contact_21_78
timestamp 1683767628
transform 1 0 15880 0 1 494
box 0 0 1 1
use contact_21  contact_21_79
timestamp 1683767628
transform 1 0 15256 0 1 370
box 0 0 1 1
use contact_21  contact_21_80
timestamp 1683767628
transform 1 0 19378 0 1 92
box 0 0 1 1
use contact_21  contact_21_81
timestamp 1683767628
transform 1 0 19842 0 1 216
box 0 0 1 1
use contact_21  contact_21_82
timestamp 1683767628
transform 1 0 19246 0 1 92
box 0 0 1 1
use contact_21  contact_21_83
timestamp 1683767628
transform 1 0 18782 0 1 216
box 0 0 1 1
use contact_21  contact_21_84
timestamp 1683767628
transform 1 0 18130 0 1 92
box 0 0 1 1
use contact_21  contact_21_85
timestamp 1683767628
transform 1 0 18594 0 1 216
box 0 0 1 1
use contact_21  contact_21_86
timestamp 1683767628
transform 1 0 17998 0 1 92
box 0 0 1 1
use contact_21  contact_21_87
timestamp 1683767628
transform 1 0 17534 0 1 216
box 0 0 1 1
use contact_21  contact_21_88
timestamp 1683767628
transform 1 0 16882 0 1 92
box 0 0 1 1
use contact_21  contact_21_89
timestamp 1683767628
transform 1 0 17346 0 1 216
box 0 0 1 1
use contact_21  contact_21_90
timestamp 1683767628
transform 1 0 16750 0 1 92
box 0 0 1 1
use contact_21  contact_21_91
timestamp 1683767628
transform 1 0 16286 0 1 216
box 0 0 1 1
use contact_21  contact_21_92
timestamp 1683767628
transform 1 0 15634 0 1 92
box 0 0 1 1
use contact_21  contact_21_93
timestamp 1683767628
transform 1 0 16098 0 1 216
box 0 0 1 1
use contact_21  contact_21_94
timestamp 1683767628
transform 1 0 15502 0 1 92
box 0 0 1 1
use contact_21  contact_21_95
timestamp 1683767628
transform 1 0 15038 0 1 216
box 0 0 1 1
use contact_21  contact_21_96
timestamp 1683767628
transform 1 0 24370 0 1 92
box 0 0 1 1
use contact_21  contact_21_97
timestamp 1683767628
transform 1 0 24834 0 1 216
box 0 0 1 1
use contact_21  contact_21_98
timestamp 1683767628
transform 1 0 24238 0 1 92
box 0 0 1 1
use contact_21  contact_21_99
timestamp 1683767628
transform 1 0 23774 0 1 216
box 0 0 1 1
use contact_21  contact_21_100
timestamp 1683767628
transform 1 0 23122 0 1 92
box 0 0 1 1
use contact_21  contact_21_101
timestamp 1683767628
transform 1 0 23586 0 1 216
box 0 0 1 1
use contact_21  contact_21_102
timestamp 1683767628
transform 1 0 22990 0 1 92
box 0 0 1 1
use contact_21  contact_21_103
timestamp 1683767628
transform 1 0 22526 0 1 216
box 0 0 1 1
use contact_21  contact_21_104
timestamp 1683767628
transform 1 0 21874 0 1 92
box 0 0 1 1
use contact_21  contact_21_105
timestamp 1683767628
transform 1 0 22338 0 1 216
box 0 0 1 1
use contact_21  contact_21_106
timestamp 1683767628
transform 1 0 21742 0 1 92
box 0 0 1 1
use contact_21  contact_21_107
timestamp 1683767628
transform 1 0 21278 0 1 216
box 0 0 1 1
use contact_21  contact_21_108
timestamp 1683767628
transform 1 0 20626 0 1 92
box 0 0 1 1
use contact_21  contact_21_109
timestamp 1683767628
transform 1 0 21090 0 1 216
box 0 0 1 1
use contact_21  contact_21_110
timestamp 1683767628
transform 1 0 20494 0 1 92
box 0 0 1 1
use contact_21  contact_21_111
timestamp 1683767628
transform 1 0 20030 0 1 216
box 0 0 1 1
use contact_21  contact_21_112
timestamp 1683767628
transform 1 0 24616 0 1 494
box 0 0 1 1
use contact_21  contact_21_113
timestamp 1683767628
transform 1 0 20872 0 1 494
box 0 0 1 1
use contact_21  contact_21_114
timestamp 1683767628
transform 1 0 23992 0 1 370
box 0 0 1 1
use contact_21  contact_21_115
timestamp 1683767628
transform 1 0 23368 0 1 494
box 0 0 1 1
use contact_21  contact_21_116
timestamp 1683767628
transform 1 0 22744 0 1 370
box 0 0 1 1
use contact_21  contact_21_117
timestamp 1683767628
transform 1 0 22120 0 1 494
box 0 0 1 1
use contact_21  contact_21_118
timestamp 1683767628
transform 1 0 21496 0 1 370
box 0 0 1 1
use contact_21  contact_21_119
timestamp 1683767628
transform 1 0 20248 0 1 370
box 0 0 1 1
use contact_21  contact_21_120
timestamp 1683767628
transform 1 0 29608 0 1 494
box 0 0 1 1
use contact_21  contact_21_121
timestamp 1683767628
transform 1 0 28984 0 1 370
box 0 0 1 1
use contact_21  contact_21_122
timestamp 1683767628
transform 1 0 28360 0 1 494
box 0 0 1 1
use contact_21  contact_21_123
timestamp 1683767628
transform 1 0 27736 0 1 370
box 0 0 1 1
use contact_21  contact_21_124
timestamp 1683767628
transform 1 0 27112 0 1 494
box 0 0 1 1
use contact_21  contact_21_125
timestamp 1683767628
transform 1 0 26488 0 1 370
box 0 0 1 1
use contact_21  contact_21_126
timestamp 1683767628
transform 1 0 25864 0 1 494
box 0 0 1 1
use contact_21  contact_21_127
timestamp 1683767628
transform 1 0 25240 0 1 370
box 0 0 1 1
use contact_21  contact_21_128
timestamp 1683767628
transform 1 0 29362 0 1 92
box 0 0 1 1
use contact_21  contact_21_129
timestamp 1683767628
transform 1 0 29826 0 1 216
box 0 0 1 1
use contact_21  contact_21_130
timestamp 1683767628
transform 1 0 29230 0 1 92
box 0 0 1 1
use contact_21  contact_21_131
timestamp 1683767628
transform 1 0 28766 0 1 216
box 0 0 1 1
use contact_21  contact_21_132
timestamp 1683767628
transform 1 0 28114 0 1 92
box 0 0 1 1
use contact_21  contact_21_133
timestamp 1683767628
transform 1 0 28578 0 1 216
box 0 0 1 1
use contact_21  contact_21_134
timestamp 1683767628
transform 1 0 27982 0 1 92
box 0 0 1 1
use contact_21  contact_21_135
timestamp 1683767628
transform 1 0 27518 0 1 216
box 0 0 1 1
use contact_21  contact_21_136
timestamp 1683767628
transform 1 0 26866 0 1 92
box 0 0 1 1
use contact_21  contact_21_137
timestamp 1683767628
transform 1 0 27330 0 1 216
box 0 0 1 1
use contact_21  contact_21_138
timestamp 1683767628
transform 1 0 26734 0 1 92
box 0 0 1 1
use contact_21  contact_21_139
timestamp 1683767628
transform 1 0 26270 0 1 216
box 0 0 1 1
use contact_21  contact_21_140
timestamp 1683767628
transform 1 0 25618 0 1 92
box 0 0 1 1
use contact_21  contact_21_141
timestamp 1683767628
transform 1 0 26082 0 1 216
box 0 0 1 1
use contact_21  contact_21_142
timestamp 1683767628
transform 1 0 25486 0 1 92
box 0 0 1 1
use contact_21  contact_21_143
timestamp 1683767628
transform 1 0 25022 0 1 216
box 0 0 1 1
use contact_21  contact_21_144
timestamp 1683767628
transform 1 0 33352 0 1 494
box 0 0 1 1
use contact_21  contact_21_145
timestamp 1683767628
transform 1 0 32728 0 1 370
box 0 0 1 1
use contact_21  contact_21_146
timestamp 1683767628
transform 1 0 32104 0 1 494
box 0 0 1 1
use contact_21  contact_21_147
timestamp 1683767628
transform 1 0 31480 0 1 370
box 0 0 1 1
use contact_21  contact_21_148
timestamp 1683767628
transform 1 0 30232 0 1 370
box 0 0 1 1
use contact_21  contact_21_149
timestamp 1683767628
transform 1 0 34354 0 1 92
box 0 0 1 1
use contact_21  contact_21_150
timestamp 1683767628
transform 1 0 34818 0 1 216
box 0 0 1 1
use contact_21  contact_21_151
timestamp 1683767628
transform 1 0 34222 0 1 92
box 0 0 1 1
use contact_21  contact_21_152
timestamp 1683767628
transform 1 0 33758 0 1 216
box 0 0 1 1
use contact_21  contact_21_153
timestamp 1683767628
transform 1 0 33106 0 1 92
box 0 0 1 1
use contact_21  contact_21_154
timestamp 1683767628
transform 1 0 33570 0 1 216
box 0 0 1 1
use contact_21  contact_21_155
timestamp 1683767628
transform 1 0 32974 0 1 92
box 0 0 1 1
use contact_21  contact_21_156
timestamp 1683767628
transform 1 0 32510 0 1 216
box 0 0 1 1
use contact_21  contact_21_157
timestamp 1683767628
transform 1 0 31858 0 1 92
box 0 0 1 1
use contact_21  contact_21_158
timestamp 1683767628
transform 1 0 32322 0 1 216
box 0 0 1 1
use contact_21  contact_21_159
timestamp 1683767628
transform 1 0 31726 0 1 92
box 0 0 1 1
use contact_21  contact_21_160
timestamp 1683767628
transform 1 0 31262 0 1 216
box 0 0 1 1
use contact_21  contact_21_161
timestamp 1683767628
transform 1 0 30610 0 1 92
box 0 0 1 1
use contact_21  contact_21_162
timestamp 1683767628
transform 1 0 31074 0 1 216
box 0 0 1 1
use contact_21  contact_21_163
timestamp 1683767628
transform 1 0 30478 0 1 92
box 0 0 1 1
use contact_21  contact_21_164
timestamp 1683767628
transform 1 0 30014 0 1 216
box 0 0 1 1
use contact_21  contact_21_165
timestamp 1683767628
transform 1 0 34600 0 1 494
box 0 0 1 1
use contact_21  contact_21_166
timestamp 1683767628
transform 1 0 30856 0 1 494
box 0 0 1 1
use contact_21  contact_21_167
timestamp 1683767628
transform 1 0 33976 0 1 370
box 0 0 1 1
use contact_21  contact_21_168
timestamp 1683767628
transform 1 0 39346 0 1 92
box 0 0 1 1
use contact_21  contact_21_169
timestamp 1683767628
transform 1 0 39810 0 1 216
box 0 0 1 1
use contact_21  contact_21_170
timestamp 1683767628
transform 1 0 39214 0 1 92
box 0 0 1 1
use contact_21  contact_21_171
timestamp 1683767628
transform 1 0 38750 0 1 216
box 0 0 1 1
use contact_21  contact_21_172
timestamp 1683767628
transform 1 0 38098 0 1 92
box 0 0 1 1
use contact_21  contact_21_173
timestamp 1683767628
transform 1 0 38562 0 1 216
box 0 0 1 1
use contact_21  contact_21_174
timestamp 1683767628
transform 1 0 37966 0 1 92
box 0 0 1 1
use contact_21  contact_21_175
timestamp 1683767628
transform 1 0 37502 0 1 216
box 0 0 1 1
use contact_21  contact_21_176
timestamp 1683767628
transform 1 0 36850 0 1 92
box 0 0 1 1
use contact_21  contact_21_177
timestamp 1683767628
transform 1 0 37314 0 1 216
box 0 0 1 1
use contact_21  contact_21_178
timestamp 1683767628
transform 1 0 36718 0 1 92
box 0 0 1 1
use contact_21  contact_21_179
timestamp 1683767628
transform 1 0 36254 0 1 216
box 0 0 1 1
use contact_21  contact_21_180
timestamp 1683767628
transform 1 0 35602 0 1 92
box 0 0 1 1
use contact_21  contact_21_181
timestamp 1683767628
transform 1 0 36066 0 1 216
box 0 0 1 1
use contact_21  contact_21_182
timestamp 1683767628
transform 1 0 35470 0 1 92
box 0 0 1 1
use contact_21  contact_21_183
timestamp 1683767628
transform 1 0 35006 0 1 216
box 0 0 1 1
use contact_21  contact_21_184
timestamp 1683767628
transform 1 0 39592 0 1 494
box 0 0 1 1
use contact_21  contact_21_185
timestamp 1683767628
transform 1 0 38968 0 1 370
box 0 0 1 1
use contact_21  contact_21_186
timestamp 1683767628
transform 1 0 38344 0 1 494
box 0 0 1 1
use contact_21  contact_21_187
timestamp 1683767628
transform 1 0 37720 0 1 370
box 0 0 1 1
use contact_21  contact_21_188
timestamp 1683767628
transform 1 0 37096 0 1 494
box 0 0 1 1
use contact_21  contact_21_189
timestamp 1683767628
transform 1 0 36472 0 1 370
box 0 0 1 1
use contact_21  contact_21_190
timestamp 1683767628
transform 1 0 35848 0 1 494
box 0 0 1 1
use contact_21  contact_21_191
timestamp 1683767628
transform 1 0 35224 0 1 370
box 0 0 1 1
use contact_22  contact_22_0
timestamp 1683767628
transform 1 0 4023 0 1 365
box 0 0 1 1
use contact_22  contact_22_1
timestamp 1683767628
transform 1 0 2775 0 1 365
box 0 0 1 1
use contact_22  contact_22_2
timestamp 1683767628
transform 1 0 279 0 1 365
box 0 0 1 1
use contact_22  contact_22_3
timestamp 1683767628
transform 1 0 1527 0 1 365
box 0 0 1 1
use contact_22  contact_22_4
timestamp 1683767628
transform 1 0 4647 0 1 489
box 0 0 1 1
use contact_22  contact_22_5
timestamp 1683767628
transform 1 0 3399 0 1 489
box 0 0 1 1
use contact_22  contact_22_6
timestamp 1683767628
transform 1 0 2151 0 1 489
box 0 0 1 1
use contact_22  contact_22_7
timestamp 1683767628
transform 1 0 903 0 1 489
box 0 0 1 1
use contact_22  contact_22_8
timestamp 1683767628
transform 1 0 4401 0 1 87
box 0 0 1 1
use contact_22  contact_22_9
timestamp 1683767628
transform 1 0 4865 0 1 211
box 0 0 1 1
use contact_22  contact_22_10
timestamp 1683767628
transform 1 0 4269 0 1 87
box 0 0 1 1
use contact_22  contact_22_11
timestamp 1683767628
transform 1 0 3805 0 1 211
box 0 0 1 1
use contact_22  contact_22_12
timestamp 1683767628
transform 1 0 3153 0 1 87
box 0 0 1 1
use contact_22  contact_22_13
timestamp 1683767628
transform 1 0 3617 0 1 211
box 0 0 1 1
use contact_22  contact_22_14
timestamp 1683767628
transform 1 0 3021 0 1 87
box 0 0 1 1
use contact_22  contact_22_15
timestamp 1683767628
transform 1 0 2557 0 1 211
box 0 0 1 1
use contact_22  contact_22_16
timestamp 1683767628
transform 1 0 1905 0 1 87
box 0 0 1 1
use contact_22  contact_22_17
timestamp 1683767628
transform 1 0 2369 0 1 211
box 0 0 1 1
use contact_22  contact_22_18
timestamp 1683767628
transform 1 0 1773 0 1 87
box 0 0 1 1
use contact_22  contact_22_19
timestamp 1683767628
transform 1 0 1309 0 1 211
box 0 0 1 1
use contact_22  contact_22_20
timestamp 1683767628
transform 1 0 657 0 1 87
box 0 0 1 1
use contact_22  contact_22_21
timestamp 1683767628
transform 1 0 1121 0 1 211
box 0 0 1 1
use contact_22  contact_22_22
timestamp 1683767628
transform 1 0 525 0 1 87
box 0 0 1 1
use contact_22  contact_22_23
timestamp 1683767628
transform 1 0 61 0 1 211
box 0 0 1 1
use contact_22  contact_22_24
timestamp 1683767628
transform 1 0 9015 0 1 365
box 0 0 1 1
use contact_22  contact_22_25
timestamp 1683767628
transform 1 0 7767 0 1 365
box 0 0 1 1
use contact_22  contact_22_26
timestamp 1683767628
transform 1 0 6519 0 1 365
box 0 0 1 1
use contact_22  contact_22_27
timestamp 1683767628
transform 1 0 5271 0 1 365
box 0 0 1 1
use contact_22  contact_22_28
timestamp 1683767628
transform 1 0 9639 0 1 489
box 0 0 1 1
use contact_22  contact_22_29
timestamp 1683767628
transform 1 0 8391 0 1 489
box 0 0 1 1
use contact_22  contact_22_30
timestamp 1683767628
transform 1 0 7143 0 1 489
box 0 0 1 1
use contact_22  contact_22_31
timestamp 1683767628
transform 1 0 5895 0 1 489
box 0 0 1 1
use contact_22  contact_22_32
timestamp 1683767628
transform 1 0 9393 0 1 87
box 0 0 1 1
use contact_22  contact_22_33
timestamp 1683767628
transform 1 0 9857 0 1 211
box 0 0 1 1
use contact_22  contact_22_34
timestamp 1683767628
transform 1 0 9261 0 1 87
box 0 0 1 1
use contact_22  contact_22_35
timestamp 1683767628
transform 1 0 8797 0 1 211
box 0 0 1 1
use contact_22  contact_22_36
timestamp 1683767628
transform 1 0 8145 0 1 87
box 0 0 1 1
use contact_22  contact_22_37
timestamp 1683767628
transform 1 0 8609 0 1 211
box 0 0 1 1
use contact_22  contact_22_38
timestamp 1683767628
transform 1 0 8013 0 1 87
box 0 0 1 1
use contact_22  contact_22_39
timestamp 1683767628
transform 1 0 7549 0 1 211
box 0 0 1 1
use contact_22  contact_22_40
timestamp 1683767628
transform 1 0 6897 0 1 87
box 0 0 1 1
use contact_22  contact_22_41
timestamp 1683767628
transform 1 0 7361 0 1 211
box 0 0 1 1
use contact_22  contact_22_42
timestamp 1683767628
transform 1 0 6765 0 1 87
box 0 0 1 1
use contact_22  contact_22_43
timestamp 1683767628
transform 1 0 6301 0 1 211
box 0 0 1 1
use contact_22  contact_22_44
timestamp 1683767628
transform 1 0 5649 0 1 87
box 0 0 1 1
use contact_22  contact_22_45
timestamp 1683767628
transform 1 0 6113 0 1 211
box 0 0 1 1
use contact_22  contact_22_46
timestamp 1683767628
transform 1 0 5517 0 1 87
box 0 0 1 1
use contact_22  contact_22_47
timestamp 1683767628
transform 1 0 5053 0 1 211
box 0 0 1 1
use contact_22  contact_22_48
timestamp 1683767628
transform 1 0 14385 0 1 87
box 0 0 1 1
use contact_22  contact_22_49
timestamp 1683767628
transform 1 0 14849 0 1 211
box 0 0 1 1
use contact_22  contact_22_50
timestamp 1683767628
transform 1 0 14253 0 1 87
box 0 0 1 1
use contact_22  contact_22_51
timestamp 1683767628
transform 1 0 13789 0 1 211
box 0 0 1 1
use contact_22  contact_22_52
timestamp 1683767628
transform 1 0 13137 0 1 87
box 0 0 1 1
use contact_22  contact_22_53
timestamp 1683767628
transform 1 0 13601 0 1 211
box 0 0 1 1
use contact_22  contact_22_54
timestamp 1683767628
transform 1 0 13005 0 1 87
box 0 0 1 1
use contact_22  contact_22_55
timestamp 1683767628
transform 1 0 12541 0 1 211
box 0 0 1 1
use contact_22  contact_22_56
timestamp 1683767628
transform 1 0 11889 0 1 87
box 0 0 1 1
use contact_22  contact_22_57
timestamp 1683767628
transform 1 0 12353 0 1 211
box 0 0 1 1
use contact_22  contact_22_58
timestamp 1683767628
transform 1 0 11757 0 1 87
box 0 0 1 1
use contact_22  contact_22_59
timestamp 1683767628
transform 1 0 11293 0 1 211
box 0 0 1 1
use contact_22  contact_22_60
timestamp 1683767628
transform 1 0 10641 0 1 87
box 0 0 1 1
use contact_22  contact_22_61
timestamp 1683767628
transform 1 0 11105 0 1 211
box 0 0 1 1
use contact_22  contact_22_62
timestamp 1683767628
transform 1 0 10509 0 1 87
box 0 0 1 1
use contact_22  contact_22_63
timestamp 1683767628
transform 1 0 10045 0 1 211
box 0 0 1 1
use contact_22  contact_22_64
timestamp 1683767628
transform 1 0 14007 0 1 365
box 0 0 1 1
use contact_22  contact_22_65
timestamp 1683767628
transform 1 0 12759 0 1 365
box 0 0 1 1
use contact_22  contact_22_66
timestamp 1683767628
transform 1 0 10263 0 1 365
box 0 0 1 1
use contact_22  contact_22_67
timestamp 1683767628
transform 1 0 11511 0 1 365
box 0 0 1 1
use contact_22  contact_22_68
timestamp 1683767628
transform 1 0 14631 0 1 489
box 0 0 1 1
use contact_22  contact_22_69
timestamp 1683767628
transform 1 0 13383 0 1 489
box 0 0 1 1
use contact_22  contact_22_70
timestamp 1683767628
transform 1 0 12135 0 1 489
box 0 0 1 1
use contact_22  contact_22_71
timestamp 1683767628
transform 1 0 10887 0 1 489
box 0 0 1 1
use contact_22  contact_22_72
timestamp 1683767628
transform 1 0 18999 0 1 365
box 0 0 1 1
use contact_22  contact_22_73
timestamp 1683767628
transform 1 0 17751 0 1 365
box 0 0 1 1
use contact_22  contact_22_74
timestamp 1683767628
transform 1 0 16503 0 1 365
box 0 0 1 1
use contact_22  contact_22_75
timestamp 1683767628
transform 1 0 15255 0 1 365
box 0 0 1 1
use contact_22  contact_22_76
timestamp 1683767628
transform 1 0 19623 0 1 489
box 0 0 1 1
use contact_22  contact_22_77
timestamp 1683767628
transform 1 0 18375 0 1 489
box 0 0 1 1
use contact_22  contact_22_78
timestamp 1683767628
transform 1 0 17127 0 1 489
box 0 0 1 1
use contact_22  contact_22_79
timestamp 1683767628
transform 1 0 15879 0 1 489
box 0 0 1 1
use contact_22  contact_22_80
timestamp 1683767628
transform 1 0 19377 0 1 87
box 0 0 1 1
use contact_22  contact_22_81
timestamp 1683767628
transform 1 0 19841 0 1 211
box 0 0 1 1
use contact_22  contact_22_82
timestamp 1683767628
transform 1 0 19245 0 1 87
box 0 0 1 1
use contact_22  contact_22_83
timestamp 1683767628
transform 1 0 18781 0 1 211
box 0 0 1 1
use contact_22  contact_22_84
timestamp 1683767628
transform 1 0 18129 0 1 87
box 0 0 1 1
use contact_22  contact_22_85
timestamp 1683767628
transform 1 0 18593 0 1 211
box 0 0 1 1
use contact_22  contact_22_86
timestamp 1683767628
transform 1 0 17997 0 1 87
box 0 0 1 1
use contact_22  contact_22_87
timestamp 1683767628
transform 1 0 17533 0 1 211
box 0 0 1 1
use contact_22  contact_22_88
timestamp 1683767628
transform 1 0 16881 0 1 87
box 0 0 1 1
use contact_22  contact_22_89
timestamp 1683767628
transform 1 0 17345 0 1 211
box 0 0 1 1
use contact_22  contact_22_90
timestamp 1683767628
transform 1 0 16749 0 1 87
box 0 0 1 1
use contact_22  contact_22_91
timestamp 1683767628
transform 1 0 16285 0 1 211
box 0 0 1 1
use contact_22  contact_22_92
timestamp 1683767628
transform 1 0 15633 0 1 87
box 0 0 1 1
use contact_22  contact_22_93
timestamp 1683767628
transform 1 0 16097 0 1 211
box 0 0 1 1
use contact_22  contact_22_94
timestamp 1683767628
transform 1 0 15501 0 1 87
box 0 0 1 1
use contact_22  contact_22_95
timestamp 1683767628
transform 1 0 15037 0 1 211
box 0 0 1 1
use contact_22  contact_22_96
timestamp 1683767628
transform 1 0 24369 0 1 87
box 0 0 1 1
use contact_22  contact_22_97
timestamp 1683767628
transform 1 0 24833 0 1 211
box 0 0 1 1
use contact_22  contact_22_98
timestamp 1683767628
transform 1 0 24237 0 1 87
box 0 0 1 1
use contact_22  contact_22_99
timestamp 1683767628
transform 1 0 23773 0 1 211
box 0 0 1 1
use contact_22  contact_22_100
timestamp 1683767628
transform 1 0 23121 0 1 87
box 0 0 1 1
use contact_22  contact_22_101
timestamp 1683767628
transform 1 0 23585 0 1 211
box 0 0 1 1
use contact_22  contact_22_102
timestamp 1683767628
transform 1 0 22989 0 1 87
box 0 0 1 1
use contact_22  contact_22_103
timestamp 1683767628
transform 1 0 22525 0 1 211
box 0 0 1 1
use contact_22  contact_22_104
timestamp 1683767628
transform 1 0 21873 0 1 87
box 0 0 1 1
use contact_22  contact_22_105
timestamp 1683767628
transform 1 0 22337 0 1 211
box 0 0 1 1
use contact_22  contact_22_106
timestamp 1683767628
transform 1 0 21741 0 1 87
box 0 0 1 1
use contact_22  contact_22_107
timestamp 1683767628
transform 1 0 21277 0 1 211
box 0 0 1 1
use contact_22  contact_22_108
timestamp 1683767628
transform 1 0 20625 0 1 87
box 0 0 1 1
use contact_22  contact_22_109
timestamp 1683767628
transform 1 0 21089 0 1 211
box 0 0 1 1
use contact_22  contact_22_110
timestamp 1683767628
transform 1 0 20493 0 1 87
box 0 0 1 1
use contact_22  contact_22_111
timestamp 1683767628
transform 1 0 20029 0 1 211
box 0 0 1 1
use contact_22  contact_22_112
timestamp 1683767628
transform 1 0 23991 0 1 365
box 0 0 1 1
use contact_22  contact_22_113
timestamp 1683767628
transform 1 0 22743 0 1 365
box 0 0 1 1
use contact_22  contact_22_114
timestamp 1683767628
transform 1 0 20247 0 1 365
box 0 0 1 1
use contact_22  contact_22_115
timestamp 1683767628
transform 1 0 21495 0 1 365
box 0 0 1 1
use contact_22  contact_22_116
timestamp 1683767628
transform 1 0 24615 0 1 489
box 0 0 1 1
use contact_22  contact_22_117
timestamp 1683767628
transform 1 0 23367 0 1 489
box 0 0 1 1
use contact_22  contact_22_118
timestamp 1683767628
transform 1 0 22119 0 1 489
box 0 0 1 1
use contact_22  contact_22_119
timestamp 1683767628
transform 1 0 20871 0 1 489
box 0 0 1 1
use contact_22  contact_22_120
timestamp 1683767628
transform 1 0 28983 0 1 365
box 0 0 1 1
use contact_22  contact_22_121
timestamp 1683767628
transform 1 0 27735 0 1 365
box 0 0 1 1
use contact_22  contact_22_122
timestamp 1683767628
transform 1 0 26487 0 1 365
box 0 0 1 1
use contact_22  contact_22_123
timestamp 1683767628
transform 1 0 25239 0 1 365
box 0 0 1 1
use contact_22  contact_22_124
timestamp 1683767628
transform 1 0 29607 0 1 489
box 0 0 1 1
use contact_22  contact_22_125
timestamp 1683767628
transform 1 0 28359 0 1 489
box 0 0 1 1
use contact_22  contact_22_126
timestamp 1683767628
transform 1 0 27111 0 1 489
box 0 0 1 1
use contact_22  contact_22_127
timestamp 1683767628
transform 1 0 25863 0 1 489
box 0 0 1 1
use contact_22  contact_22_128
timestamp 1683767628
transform 1 0 29361 0 1 87
box 0 0 1 1
use contact_22  contact_22_129
timestamp 1683767628
transform 1 0 29825 0 1 211
box 0 0 1 1
use contact_22  contact_22_130
timestamp 1683767628
transform 1 0 29229 0 1 87
box 0 0 1 1
use contact_22  contact_22_131
timestamp 1683767628
transform 1 0 28765 0 1 211
box 0 0 1 1
use contact_22  contact_22_132
timestamp 1683767628
transform 1 0 28113 0 1 87
box 0 0 1 1
use contact_22  contact_22_133
timestamp 1683767628
transform 1 0 28577 0 1 211
box 0 0 1 1
use contact_22  contact_22_134
timestamp 1683767628
transform 1 0 27981 0 1 87
box 0 0 1 1
use contact_22  contact_22_135
timestamp 1683767628
transform 1 0 27517 0 1 211
box 0 0 1 1
use contact_22  contact_22_136
timestamp 1683767628
transform 1 0 26865 0 1 87
box 0 0 1 1
use contact_22  contact_22_137
timestamp 1683767628
transform 1 0 27329 0 1 211
box 0 0 1 1
use contact_22  contact_22_138
timestamp 1683767628
transform 1 0 26733 0 1 87
box 0 0 1 1
use contact_22  contact_22_139
timestamp 1683767628
transform 1 0 26269 0 1 211
box 0 0 1 1
use contact_22  contact_22_140
timestamp 1683767628
transform 1 0 25617 0 1 87
box 0 0 1 1
use contact_22  contact_22_141
timestamp 1683767628
transform 1 0 26081 0 1 211
box 0 0 1 1
use contact_22  contact_22_142
timestamp 1683767628
transform 1 0 25485 0 1 87
box 0 0 1 1
use contact_22  contact_22_143
timestamp 1683767628
transform 1 0 25021 0 1 211
box 0 0 1 1
use contact_22  contact_22_144
timestamp 1683767628
transform 1 0 32727 0 1 365
box 0 0 1 1
use contact_22  contact_22_145
timestamp 1683767628
transform 1 0 30231 0 1 365
box 0 0 1 1
use contact_22  contact_22_146
timestamp 1683767628
transform 1 0 31479 0 1 365
box 0 0 1 1
use contact_22  contact_22_147
timestamp 1683767628
transform 1 0 34599 0 1 489
box 0 0 1 1
use contact_22  contact_22_148
timestamp 1683767628
transform 1 0 33351 0 1 489
box 0 0 1 1
use contact_22  contact_22_149
timestamp 1683767628
transform 1 0 32103 0 1 489
box 0 0 1 1
use contact_22  contact_22_150
timestamp 1683767628
transform 1 0 30855 0 1 489
box 0 0 1 1
use contact_22  contact_22_151
timestamp 1683767628
transform 1 0 34353 0 1 87
box 0 0 1 1
use contact_22  contact_22_152
timestamp 1683767628
transform 1 0 34817 0 1 211
box 0 0 1 1
use contact_22  contact_22_153
timestamp 1683767628
transform 1 0 34221 0 1 87
box 0 0 1 1
use contact_22  contact_22_154
timestamp 1683767628
transform 1 0 33757 0 1 211
box 0 0 1 1
use contact_22  contact_22_155
timestamp 1683767628
transform 1 0 33105 0 1 87
box 0 0 1 1
use contact_22  contact_22_156
timestamp 1683767628
transform 1 0 33569 0 1 211
box 0 0 1 1
use contact_22  contact_22_157
timestamp 1683767628
transform 1 0 32973 0 1 87
box 0 0 1 1
use contact_22  contact_22_158
timestamp 1683767628
transform 1 0 32509 0 1 211
box 0 0 1 1
use contact_22  contact_22_159
timestamp 1683767628
transform 1 0 31857 0 1 87
box 0 0 1 1
use contact_22  contact_22_160
timestamp 1683767628
transform 1 0 32321 0 1 211
box 0 0 1 1
use contact_22  contact_22_161
timestamp 1683767628
transform 1 0 31725 0 1 87
box 0 0 1 1
use contact_22  contact_22_162
timestamp 1683767628
transform 1 0 31261 0 1 211
box 0 0 1 1
use contact_22  contact_22_163
timestamp 1683767628
transform 1 0 30609 0 1 87
box 0 0 1 1
use contact_22  contact_22_164
timestamp 1683767628
transform 1 0 31073 0 1 211
box 0 0 1 1
use contact_22  contact_22_165
timestamp 1683767628
transform 1 0 30477 0 1 87
box 0 0 1 1
use contact_22  contact_22_166
timestamp 1683767628
transform 1 0 30013 0 1 211
box 0 0 1 1
use contact_22  contact_22_167
timestamp 1683767628
transform 1 0 33975 0 1 365
box 0 0 1 1
use contact_22  contact_22_168
timestamp 1683767628
transform 1 0 39345 0 1 87
box 0 0 1 1
use contact_22  contact_22_169
timestamp 1683767628
transform 1 0 39809 0 1 211
box 0 0 1 1
use contact_22  contact_22_170
timestamp 1683767628
transform 1 0 39213 0 1 87
box 0 0 1 1
use contact_22  contact_22_171
timestamp 1683767628
transform 1 0 38749 0 1 211
box 0 0 1 1
use contact_22  contact_22_172
timestamp 1683767628
transform 1 0 38097 0 1 87
box 0 0 1 1
use contact_22  contact_22_173
timestamp 1683767628
transform 1 0 38561 0 1 211
box 0 0 1 1
use contact_22  contact_22_174
timestamp 1683767628
transform 1 0 37965 0 1 87
box 0 0 1 1
use contact_22  contact_22_175
timestamp 1683767628
transform 1 0 37501 0 1 211
box 0 0 1 1
use contact_22  contact_22_176
timestamp 1683767628
transform 1 0 36849 0 1 87
box 0 0 1 1
use contact_22  contact_22_177
timestamp 1683767628
transform 1 0 37313 0 1 211
box 0 0 1 1
use contact_22  contact_22_178
timestamp 1683767628
transform 1 0 36717 0 1 87
box 0 0 1 1
use contact_22  contact_22_179
timestamp 1683767628
transform 1 0 36253 0 1 211
box 0 0 1 1
use contact_22  contact_22_180
timestamp 1683767628
transform 1 0 35601 0 1 87
box 0 0 1 1
use contact_22  contact_22_181
timestamp 1683767628
transform 1 0 36065 0 1 211
box 0 0 1 1
use contact_22  contact_22_182
timestamp 1683767628
transform 1 0 35469 0 1 87
box 0 0 1 1
use contact_22  contact_22_183
timestamp 1683767628
transform 1 0 35005 0 1 211
box 0 0 1 1
use contact_22  contact_22_184
timestamp 1683767628
transform 1 0 38967 0 1 365
box 0 0 1 1
use contact_22  contact_22_185
timestamp 1683767628
transform 1 0 37719 0 1 365
box 0 0 1 1
use contact_22  contact_22_186
timestamp 1683767628
transform 1 0 36471 0 1 365
box 0 0 1 1
use contact_22  contact_22_187
timestamp 1683767628
transform 1 0 35223 0 1 365
box 0 0 1 1
use contact_22  contact_22_188
timestamp 1683767628
transform 1 0 39591 0 1 489
box 0 0 1 1
use contact_22  contact_22_189
timestamp 1683767628
transform 1 0 38343 0 1 489
box 0 0 1 1
use contact_22  contact_22_190
timestamp 1683767628
transform 1 0 37095 0 1 489
box 0 0 1 1
use contact_22  contact_22_191
timestamp 1683767628
transform 1 0 35847 0 1 489
box 0 0 1 1
use single_level_column_mux  single_level_column_mux_0
timestamp 1683767628
transform -1 0 4992 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_1
timestamp 1683767628
transform 1 0 3744 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_2
timestamp 1683767628
transform -1 0 3744 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_3
timestamp 1683767628
transform 1 0 2496 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_4
timestamp 1683767628
transform -1 0 2496 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_5
timestamp 1683767628
transform 1 0 1248 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_6
timestamp 1683767628
transform -1 0 1248 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_7
timestamp 1683767628
transform 1 0 0 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_8
timestamp 1683767628
transform -1 0 9984 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_9
timestamp 1683767628
transform 1 0 8736 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_10
timestamp 1683767628
transform -1 0 8736 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_11
timestamp 1683767628
transform 1 0 7488 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_12
timestamp 1683767628
transform -1 0 7488 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_13
timestamp 1683767628
transform 1 0 6240 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_14
timestamp 1683767628
transform -1 0 6240 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_15
timestamp 1683767628
transform 1 0 4992 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_16
timestamp 1683767628
transform -1 0 14976 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_17
timestamp 1683767628
transform 1 0 13728 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_18
timestamp 1683767628
transform -1 0 13728 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_19
timestamp 1683767628
transform 1 0 12480 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_20
timestamp 1683767628
transform -1 0 12480 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_21
timestamp 1683767628
transform 1 0 11232 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_22
timestamp 1683767628
transform -1 0 11232 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_23
timestamp 1683767628
transform 1 0 9984 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_24
timestamp 1683767628
transform -1 0 19968 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_25
timestamp 1683767628
transform 1 0 18720 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_26
timestamp 1683767628
transform -1 0 18720 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_27
timestamp 1683767628
transform 1 0 17472 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_28
timestamp 1683767628
transform -1 0 17472 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_29
timestamp 1683767628
transform 1 0 16224 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_30
timestamp 1683767628
transform -1 0 16224 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_31
timestamp 1683767628
transform 1 0 14976 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_32
timestamp 1683767628
transform -1 0 24960 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_33
timestamp 1683767628
transform 1 0 23712 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_34
timestamp 1683767628
transform -1 0 23712 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_35
timestamp 1683767628
transform 1 0 22464 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_36
timestamp 1683767628
transform -1 0 22464 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_37
timestamp 1683767628
transform 1 0 21216 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_38
timestamp 1683767628
transform -1 0 21216 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_39
timestamp 1683767628
transform 1 0 19968 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_40
timestamp 1683767628
transform -1 0 29952 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_41
timestamp 1683767628
transform 1 0 28704 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_42
timestamp 1683767628
transform -1 0 28704 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_43
timestamp 1683767628
transform 1 0 27456 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_44
timestamp 1683767628
transform -1 0 27456 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_45
timestamp 1683767628
transform 1 0 26208 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_46
timestamp 1683767628
transform -1 0 26208 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_47
timestamp 1683767628
transform 1 0 24960 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_48
timestamp 1683767628
transform -1 0 34944 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_49
timestamp 1683767628
transform 1 0 33696 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_50
timestamp 1683767628
transform -1 0 33696 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_51
timestamp 1683767628
transform 1 0 32448 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_52
timestamp 1683767628
transform -1 0 32448 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_53
timestamp 1683767628
transform 1 0 31200 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_54
timestamp 1683767628
transform -1 0 31200 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_55
timestamp 1683767628
transform 1 0 29952 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_56
timestamp 1683767628
transform -1 0 39936 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_57
timestamp 1683767628
transform 1 0 38688 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_58
timestamp 1683767628
transform -1 0 38688 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_59
timestamp 1683767628
transform 1 0 37440 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_60
timestamp 1683767628
transform -1 0 37440 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_61
timestamp 1683767628
transform 1 0 36192 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_62
timestamp 1683767628
transform -1 0 36192 0 1 620
box 65 0 675 1364
use single_level_column_mux  single_level_column_mux_63
timestamp 1683767628
transform 1 0 34944 0 1 620
box 65 0 675 1364
<< labels >>
rlabel metal1 s 27550 1956 27550 1956 4 bl_44
port 89 nsew
rlabel metal1 s 29262 1956 29262 1956 4 br_46
port 94 nsew
rlabel metal1 s 21906 1956 21906 1956 4 br_35
port 72 nsew
rlabel metal1 s 34254 1956 34254 1956 4 br_54
port 110 nsew
rlabel metal1 s 28146 1956 28146 1956 4 br_45
port 92 nsew
rlabel metal1 s 34386 1956 34386 1956 4 br_55
port 112 nsew
rlabel metal1 s 36098 1956 36098 1956 4 bl_57
port 115 nsew
rlabel metal1 s 35634 1956 35634 1956 4 br_57
port 116 nsew
rlabel metal1 s 38782 1956 38782 1956 4 bl_62
port 125 nsew
rlabel metal1 s 21310 1956 21310 1956 4 bl_34
port 69 nsew
rlabel metal1 s 35038 1956 35038 1956 4 bl_56
port 113 nsew
rlabel metal1 s 29858 1956 29858 1956 4 bl_47
port 95 nsew
rlabel metal1 s 37346 1956 37346 1956 4 bl_59
port 119 nsew
rlabel metal1 s 39842 1956 39842 1956 4 bl_63
port 127 nsew
rlabel metal1 s 26302 1956 26302 1956 4 bl_42
port 85 nsew
rlabel metal1 s 33006 1956 33006 1956 4 br_52
port 106 nsew
rlabel metal1 s 32542 1956 32542 1956 4 bl_52
port 105 nsew
rlabel metal1 s 34850 1956 34850 1956 4 bl_55
port 111 nsew
rlabel metal1 s 22370 1956 22370 1956 4 bl_35
port 71 nsew
rlabel metal1 s 30046 1956 30046 1956 4 bl_48
port 97 nsew
rlabel metal1 s 25518 1956 25518 1956 4 br_40
port 82 nsew
rlabel metal1 s 23806 1956 23806 1956 4 bl_38
port 77 nsew
rlabel metal1 s 33790 1956 33790 1956 4 bl_54
port 109 nsew
rlabel metal1 s 31294 1956 31294 1956 4 bl_50
port 101 nsew
rlabel metal1 s 25054 1956 25054 1956 4 bl_40
port 81 nsew
rlabel metal1 s 24402 1956 24402 1956 4 br_39
port 80 nsew
rlabel metal1 s 26114 1956 26114 1956 4 bl_41
port 83 nsew
rlabel metal1 s 38130 1956 38130 1956 4 br_61
port 124 nsew
rlabel metal1 s 30510 1956 30510 1956 4 br_48
port 98 nsew
rlabel metal1 s 38594 1956 38594 1956 4 bl_61
port 123 nsew
rlabel metal1 s 28610 1956 28610 1956 4 bl_45
port 91 nsew
rlabel metal1 s 33602 1956 33602 1956 4 bl_53
port 107 nsew
rlabel metal1 s 20062 1956 20062 1956 4 bl_32
port 65 nsew
rlabel metal1 s 28798 1956 28798 1956 4 bl_46
port 93 nsew
rlabel metal1 s 36882 1956 36882 1956 4 br_59
port 120 nsew
rlabel metal1 s 22558 1956 22558 1956 4 bl_36
port 73 nsew
rlabel metal1 s 37998 1956 37998 1956 4 br_60
port 122 nsew
rlabel metal1 s 30642 1956 30642 1956 4 br_49
port 100 nsew
rlabel metal1 s 24866 1956 24866 1956 4 bl_39
port 79 nsew
rlabel metal1 s 23022 1956 23022 1956 4 br_36
port 74 nsew
rlabel metal1 s 37534 1956 37534 1956 4 bl_60
port 121 nsew
rlabel metal1 s 31106 1956 31106 1956 4 bl_49
port 99 nsew
rlabel metal1 s 39246 1956 39246 1956 4 br_62
port 126 nsew
rlabel metal1 s 25650 1956 25650 1956 4 br_41
port 84 nsew
rlabel metal1 s 26898 1956 26898 1956 4 br_43
port 88 nsew
rlabel metal1 s 35502 1956 35502 1956 4 br_56
port 114 nsew
rlabel metal1 s 23618 1956 23618 1956 4 bl_37
port 75 nsew
rlabel metal1 s 23154 1956 23154 1956 4 br_37
port 76 nsew
rlabel metal1 s 28014 1956 28014 1956 4 br_44
port 90 nsew
rlabel metal1 s 31890 1956 31890 1956 4 br_51
port 104 nsew
rlabel metal1 s 33138 1956 33138 1956 4 br_53
port 108 nsew
rlabel metal1 s 36750 1956 36750 1956 4 br_58
port 118 nsew
rlabel metal1 s 24270 1956 24270 1956 4 br_38
port 78 nsew
rlabel metal1 s 26766 1956 26766 1956 4 br_42
port 86 nsew
rlabel metal1 s 20526 1956 20526 1956 4 br_32
port 66 nsew
rlabel metal1 s 39378 1956 39378 1956 4 br_63
port 128 nsew
rlabel metal1 s 29394 1956 29394 1956 4 br_47
port 96 nsew
rlabel metal1 s 21122 1956 21122 1956 4 bl_33
port 67 nsew
rlabel metal1 s 21774 1956 21774 1956 4 br_34
port 70 nsew
rlabel metal1 s 27362 1956 27362 1956 4 bl_43
port 87 nsew
rlabel metal1 s 20658 1956 20658 1956 4 br_33
port 68 nsew
rlabel metal1 s 36286 1956 36286 1956 4 bl_58
port 117 nsew
rlabel metal1 s 32354 1956 32354 1956 4 bl_51
port 103 nsew
rlabel metal1 s 31758 1956 31758 1956 4 br_50
port 102 nsew
rlabel metal1 s 25054 434 25054 434 4 bl_out_20
port 171 nsew
rlabel metal1 s 35038 434 35038 434 4 bl_out_28
port 187 nsew
rlabel metal1 s 33790 434 33790 434 4 bl_out_27
port 185 nsew
rlabel metal1 s 38782 434 38782 434 4 bl_out_31
port 193 nsew
rlabel metal1 s 23806 434 23806 434 4 bl_out_19
port 169 nsew
rlabel metal1 s 27550 434 27550 434 4 bl_out_22
port 175 nsew
rlabel metal1 s 26302 434 26302 434 4 bl_out_21
port 173 nsew
rlabel metal1 s 21310 434 21310 434 4 bl_out_17
port 165 nsew
rlabel metal1 s 37534 434 37534 434 4 bl_out_30
port 191 nsew
rlabel metal1 s 20062 434 20062 434 4 bl_out_16
port 163 nsew
rlabel metal1 s 36286 434 36286 434 4 bl_out_29
port 189 nsew
rlabel metal1 s 31294 434 31294 434 4 bl_out_25
port 181 nsew
rlabel metal1 s 32542 434 32542 434 4 bl_out_26
port 183 nsew
rlabel metal1 s 30046 434 30046 434 4 bl_out_24
port 179 nsew
rlabel metal1 s 22558 434 22558 434 4 bl_out_18
port 167 nsew
rlabel metal1 s 28798 434 28798 434 4 bl_out_23
port 177 nsew
rlabel metal1 s 7582 1956 7582 1956 4 bl_12
port 25 nsew
rlabel metal1 s 7394 1956 7394 1956 4 bl_11
port 23 nsew
rlabel metal1 s 8178 1956 8178 1956 4 br_13
port 28 nsew
rlabel metal1 s 16318 1956 16318 1956 4 bl_26
port 53 nsew
rlabel metal1 s 17378 1956 17378 1956 4 bl_27
port 55 nsew
rlabel metal1 s 10542 1956 10542 1956 4 br_16
port 34 nsew
rlabel metal1 s 1938 1956 1938 1956 4 br_3
port 8 nsew
rlabel metal1 s 10674 1956 10674 1956 4 br_17
port 36 nsew
rlabel metal1 s 19410 1956 19410 1956 4 br_31
port 64 nsew
rlabel metal1 s 2402 1956 2402 1956 4 bl_3
port 7 nsew
rlabel metal1 s 4898 1956 4898 1956 4 bl_7
port 15 nsew
rlabel metal1 s 13170 1956 13170 1956 4 br_21
port 44 nsew
rlabel metal1 s 16782 1956 16782 1956 4 br_26
port 54 nsew
rlabel metal1 s 4302 1956 4302 1956 4 br_6
port 14 nsew
rlabel metal1 s 3054 1956 3054 1956 4 br_4
port 10 nsew
rlabel metal1 s 15666 1956 15666 1956 4 br_25
port 52 nsew
rlabel metal1 s 690 1956 690 1956 4 br_1
port 4 nsew
rlabel metal1 s 18030 1956 18030 1956 4 br_28
port 58 nsew
rlabel metal1 s 5550 1956 5550 1956 4 br_8
port 18 nsew
rlabel metal1 s 18626 1956 18626 1956 4 bl_29
port 59 nsew
rlabel metal1 s 15070 1956 15070 1956 4 bl_24
port 49 nsew
rlabel metal1 s 6334 1956 6334 1956 4 bl_10
port 21 nsew
rlabel metal1 s 19278 1956 19278 1956 4 br_30
port 62 nsew
rlabel metal1 s 3650 1956 3650 1956 4 bl_5
port 11 nsew
rlabel metal1 s 5682 1956 5682 1956 4 br_9
port 20 nsew
rlabel metal1 s 13822 1956 13822 1956 4 bl_22
port 45 nsew
rlabel metal1 s 16130 1956 16130 1956 4 bl_25
port 51 nsew
rlabel metal1 s 9294 1956 9294 1956 4 br_14
port 30 nsew
rlabel metal1 s 1806 1956 1806 1956 4 br_2
port 6 nsew
rlabel metal1 s 9890 1956 9890 1956 4 bl_15
port 31 nsew
rlabel metal1 s 9426 1956 9426 1956 4 br_15
port 32 nsew
rlabel metal1 s 16914 1956 16914 1956 4 br_27
port 56 nsew
rlabel metal1 s 11922 1956 11922 1956 4 br_19
port 40 nsew
rlabel metal1 s 6146 1956 6146 1956 4 bl_9
port 19 nsew
rlabel metal1 s 14286 1956 14286 1956 4 br_22
port 46 nsew
rlabel metal1 s 8642 1956 8642 1956 4 bl_13
port 27 nsew
rlabel metal1 s 3838 1956 3838 1956 4 bl_6
port 13 nsew
rlabel metal1 s 8830 1956 8830 1956 4 bl_14
port 29 nsew
rlabel metal1 s 18162 1956 18162 1956 4 br_29
port 60 nsew
rlabel metal1 s 12574 1956 12574 1956 4 bl_20
port 41 nsew
rlabel metal1 s 558 1956 558 1956 4 br_0
port 2 nsew
rlabel metal1 s 15534 1956 15534 1956 4 br_24
port 50 nsew
rlabel metal1 s 2590 1956 2590 1956 4 bl_4
port 9 nsew
rlabel metal1 s 94 1956 94 1956 4 bl_0
port 1 nsew
rlabel metal1 s 11790 1956 11790 1956 4 br_18
port 38 nsew
rlabel metal1 s 17566 1956 17566 1956 4 bl_28
port 57 nsew
rlabel metal1 s 10078 1956 10078 1956 4 bl_16
port 33 nsew
rlabel metal1 s 14882 1956 14882 1956 4 bl_23
port 47 nsew
rlabel metal1 s 3838 434 3838 434 4 bl_out_3
port 137 nsew
rlabel metal1 s 16318 434 16318 434 4 bl_out_13
port 157 nsew
rlabel metal1 s 7582 434 7582 434 4 bl_out_6
port 143 nsew
rlabel metal1 s 2590 434 2590 434 4 bl_out_2
port 135 nsew
rlabel metal1 s 1342 434 1342 434 4 bl_out_1
port 133 nsew
rlabel metal1 s 10078 434 10078 434 4 bl_out_8
port 147 nsew
rlabel metal1 s 5086 434 5086 434 4 bl_out_4
port 139 nsew
rlabel metal1 s 12574 434 12574 434 4 bl_out_10
port 151 nsew
rlabel metal1 s 8830 434 8830 434 4 bl_out_7
port 145 nsew
rlabel metal1 s 15070 434 15070 434 4 bl_out_12
port 155 nsew
rlabel metal1 s 13822 434 13822 434 4 bl_out_11
port 153 nsew
rlabel metal1 s 6334 434 6334 434 4 bl_out_5
port 141 nsew
rlabel metal1 s 11326 434 11326 434 4 bl_out_9
port 149 nsew
rlabel metal1 s 18814 434 18814 434 4 bl_out_15
port 161 nsew
rlabel metal1 s 94 434 94 434 4 bl_out_0
port 131 nsew
rlabel metal1 s 17566 434 17566 434 4 bl_out_14
port 159 nsew
rlabel metal1 s 6930 1956 6930 1956 4 br_11
port 24 nsew
rlabel metal1 s 6798 1956 6798 1956 4 br_10
port 22 nsew
rlabel metal1 s 1342 1956 1342 1956 4 bl_2
port 5 nsew
rlabel metal1 s 8046 1956 8046 1956 4 br_12
port 26 nsew
rlabel metal1 s 5086 1956 5086 1956 4 bl_8
port 17 nsew
rlabel metal1 s 3186 1956 3186 1956 4 br_5
port 12 nsew
rlabel metal1 s 14418 1956 14418 1956 4 br_23
port 48 nsew
rlabel metal1 s 12386 1956 12386 1956 4 bl_19
port 39 nsew
rlabel metal1 s 13634 1956 13634 1956 4 bl_21
port 43 nsew
rlabel metal1 s 13038 1956 13038 1956 4 br_20
port 42 nsew
rlabel metal1 s 1154 1956 1154 1956 4 bl_1
port 3 nsew
rlabel metal1 s 4434 1956 4434 1956 4 br_7
port 16 nsew
rlabel metal1 s 18814 1956 18814 1956 4 bl_30
port 61 nsew
rlabel metal1 s 19874 1956 19874 1956 4 bl_31
port 63 nsew
rlabel metal1 s 11138 1956 11138 1956 4 bl_17
port 35 nsew
rlabel metal1 s 11326 1956 11326 1956 4 bl_18
port 37 nsew
rlabel metal1 s 1806 372 1806 372 4 br_out_1
port 134 nsew
rlabel metal1 s 11790 372 11790 372 4 br_out_9
port 150 nsew
rlabel metal1 s 6798 372 6798 372 4 br_out_5
port 142 nsew
rlabel metal1 s 10542 372 10542 372 4 br_out_8
port 148 nsew
rlabel metal1 s 4302 372 4302 372 4 br_out_3
port 138 nsew
rlabel metal1 s 3054 372 3054 372 4 br_out_2
port 136 nsew
rlabel metal1 s 18030 372 18030 372 4 br_out_14
port 160 nsew
rlabel metal1 s 16782 372 16782 372 4 br_out_13
port 158 nsew
rlabel metal1 s 5550 372 5550 372 4 br_out_4
port 140 nsew
rlabel metal1 s 558 372 558 372 4 br_out_0
port 132 nsew
rlabel metal1 s 9294 372 9294 372 4 br_out_7
port 146 nsew
rlabel metal1 s 8046 372 8046 372 4 br_out_6
port 144 nsew
rlabel metal1 s 19278 372 19278 372 4 br_out_15
port 162 nsew
rlabel metal1 s 15534 372 15534 372 4 br_out_12
port 156 nsew
rlabel metal1 s 13038 372 13038 372 4 br_out_10
port 152 nsew
rlabel metal1 s 14286 372 14286 372 4 br_out_11
port 154 nsew
rlabel metal1 s 28014 372 28014 372 4 br_out_22
port 176 nsew
rlabel metal1 s 21774 372 21774 372 4 br_out_17
port 166 nsew
rlabel metal1 s 26766 372 26766 372 4 br_out_21
port 174 nsew
rlabel metal1 s 30510 372 30510 372 4 br_out_24
port 180 nsew
rlabel metal1 s 31758 372 31758 372 4 br_out_25
port 182 nsew
rlabel metal1 s 34254 372 34254 372 4 br_out_27
port 186 nsew
rlabel metal1 s 36750 372 36750 372 4 br_out_29
port 190 nsew
rlabel metal1 s 37998 372 37998 372 4 br_out_30
port 192 nsew
rlabel metal1 s 35502 372 35502 372 4 br_out_28
port 188 nsew
rlabel metal1 s 20526 372 20526 372 4 br_out_16
port 164 nsew
rlabel metal1 s 29262 372 29262 372 4 br_out_23
port 178 nsew
rlabel metal1 s 24270 372 24270 372 4 br_out_19
port 170 nsew
rlabel metal1 s 25518 372 25518 372 4 br_out_20
port 172 nsew
rlabel metal1 s 39246 372 39246 372 4 br_out_31
port 194 nsew
rlabel metal1 s 33006 372 33006 372 4 br_out_26
port 184 nsew
rlabel metal1 s 23022 372 23022 372 4 br_out_18
port 168 nsew
rlabel metal3 s 11856 1307 11856 1307 4 gnd
port 195 nsew
rlabel metal3 s 11856 1307 11856 1307 4 gnd
port 195 nsew
rlabel metal3 s 35568 1307 35568 1307 4 gnd
port 195 nsew
rlabel metal3 s 4368 1307 4368 1307 4 gnd
port 195 nsew
rlabel metal3 s 29328 1307 29328 1307 4 gnd
port 195 nsew
rlabel metal3 s 20592 1307 20592 1307 4 gnd
port 195 nsew
rlabel metal3 s 29328 1307 29328 1307 4 gnd
port 195 nsew
rlabel metal3 s 10608 1307 10608 1307 4 gnd
port 195 nsew
rlabel metal3 s 5616 1307 5616 1307 4 gnd
port 195 nsew
rlabel metal3 s 5616 1307 5616 1307 4 gnd
port 195 nsew
rlabel metal3 s 9360 1307 9360 1307 4 gnd
port 195 nsew
rlabel metal3 s 36816 1307 36816 1307 4 gnd
port 195 nsew
rlabel metal3 s 33072 1307 33072 1307 4 gnd
port 195 nsew
rlabel metal3 s 15600 1307 15600 1307 4 gnd
port 195 nsew
rlabel metal3 s 15600 1307 15600 1307 4 gnd
port 195 nsew
rlabel metal3 s 33072 1307 33072 1307 4 gnd
port 195 nsew
rlabel metal3 s 39312 1307 39312 1307 4 gnd
port 195 nsew
rlabel metal3 s 21840 1307 21840 1307 4 gnd
port 195 nsew
rlabel metal3 s 1872 1307 1872 1307 4 gnd
port 195 nsew
rlabel metal3 s 21840 1307 21840 1307 4 gnd
port 195 nsew
rlabel metal3 s 38064 1307 38064 1307 4 gnd
port 195 nsew
rlabel metal3 s 38064 1307 38064 1307 4 gnd
port 195 nsew
rlabel metal3 s 24336 1307 24336 1307 4 gnd
port 195 nsew
rlabel metal3 s 3120 1307 3120 1307 4 gnd
port 195 nsew
rlabel metal3 s 3120 1307 3120 1307 4 gnd
port 195 nsew
rlabel metal3 s 18096 1307 18096 1307 4 gnd
port 195 nsew
rlabel metal3 s 18096 1307 18096 1307 4 gnd
port 195 nsew
rlabel metal3 s 25584 1307 25584 1307 4 gnd
port 195 nsew
rlabel metal3 s 13104 1307 13104 1307 4 gnd
port 195 nsew
rlabel metal3 s 14352 1307 14352 1307 4 gnd
port 195 nsew
rlabel metal3 s 19344 1307 19344 1307 4 gnd
port 195 nsew
rlabel metal3 s 26832 1307 26832 1307 4 gnd
port 195 nsew
rlabel metal3 s 624 1307 624 1307 4 gnd
port 195 nsew
rlabel metal3 s 16848 1307 16848 1307 4 gnd
port 195 nsew
rlabel metal3 s 8112 1307 8112 1307 4 gnd
port 195 nsew
rlabel metal3 s 23088 1307 23088 1307 4 gnd
port 195 nsew
rlabel metal3 s 6864 1307 6864 1307 4 gnd
port 195 nsew
rlabel metal3 s 6864 1307 6864 1307 4 gnd
port 195 nsew
rlabel metal3 s 28080 1307 28080 1307 4 gnd
port 195 nsew
rlabel metal3 s 30576 1307 30576 1307 4 gnd
port 195 nsew
rlabel metal3 s 31824 1307 31824 1307 4 gnd
port 195 nsew
rlabel metal3 s 34320 1307 34320 1307 4 gnd
port 195 nsew
rlabel metal3 s 19968 402 19968 402 4 sel_0
port 129 nsew
rlabel metal3 s 19968 526 19968 526 4 sel_1
port 130 nsew
<< properties >>
string FIXED_BBOX 0 0 39936 1984
string GDS_END 3593022
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 3513806
<< end >>
