magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -66 377 3810 897
<< pwell >>
rect 1022 223 1280 233
rect 1022 217 1848 223
rect 2173 217 3740 283
rect 4 43 3740 217
rect -26 -43 3770 43
<< mvnmos >>
rect 83 107 183 191
rect 239 107 339 191
rect 381 107 481 191
rect 537 107 637 191
rect 679 107 779 191
rect 835 107 935 191
rect 1101 123 1201 207
rect 1371 113 1471 197
rect 1527 113 1627 197
rect 1669 113 1769 197
rect 1935 107 2035 191
rect 2077 107 2177 191
rect 2252 107 2352 257
rect 2394 107 2494 257
rect 2569 173 2669 257
rect 2712 173 2812 257
rect 2854 173 2954 257
rect 3043 173 3143 257
rect 3378 173 3478 257
rect 3557 107 3657 257
<< mvpmos >>
rect 83 569 183 653
rect 239 569 339 653
rect 381 569 481 653
rect 537 569 637 653
rect 679 569 779 653
rect 858 569 958 719
rect 1156 533 1256 683
rect 1430 543 1530 627
rect 1586 543 1686 627
rect 1728 543 1828 627
rect 1900 543 2000 627
rect 2056 543 2156 627
rect 2235 543 2335 743
rect 2377 543 2477 743
rect 2556 543 2656 627
rect 2698 543 2798 627
rect 2854 543 2954 627
rect 3120 613 3220 697
rect 3386 475 3486 625
rect 3561 475 3661 675
<< mvndiff >>
rect 30 166 83 191
rect 30 132 38 166
rect 72 132 83 166
rect 30 107 83 132
rect 183 166 239 191
rect 183 132 194 166
rect 228 132 239 166
rect 183 107 239 132
rect 339 107 381 191
rect 481 166 537 191
rect 481 132 492 166
rect 526 132 537 166
rect 481 107 537 132
rect 637 107 679 191
rect 779 166 835 191
rect 779 132 790 166
rect 824 132 835 166
rect 779 107 835 132
rect 935 166 988 191
rect 935 132 946 166
rect 980 132 988 166
rect 935 107 988 132
rect 1048 182 1101 207
rect 1048 148 1056 182
rect 1090 148 1101 182
rect 1048 123 1101 148
rect 1201 182 1254 207
rect 1201 148 1212 182
rect 1246 148 1254 182
rect 1201 123 1254 148
rect 1314 173 1371 197
rect 1314 139 1326 173
rect 1360 139 1371 173
rect 1314 113 1371 139
rect 1471 172 1527 197
rect 1471 138 1482 172
rect 1516 138 1527 172
rect 1471 113 1527 138
rect 1627 113 1669 197
rect 1769 172 1822 197
rect 2199 191 2252 257
rect 1769 138 1780 172
rect 1814 138 1822 172
rect 1769 113 1822 138
rect 1882 166 1935 191
rect 1882 132 1890 166
rect 1924 132 1935 166
rect 1882 107 1935 132
rect 2035 107 2077 191
rect 2177 176 2252 191
rect 2177 142 2207 176
rect 2241 142 2252 176
rect 2177 107 2252 142
rect 2352 107 2394 257
rect 2494 229 2569 257
rect 2494 195 2505 229
rect 2539 195 2569 229
rect 2494 173 2569 195
rect 2669 173 2712 257
rect 2812 173 2854 257
rect 2954 232 3043 257
rect 2954 198 2965 232
rect 2999 198 3043 232
rect 2954 173 3043 198
rect 3143 232 3200 257
rect 3143 198 3154 232
rect 3188 198 3200 232
rect 3143 173 3200 198
rect 3321 232 3378 257
rect 3321 198 3333 232
rect 3367 198 3378 232
rect 3321 173 3378 198
rect 3478 249 3557 257
rect 3478 215 3512 249
rect 3546 215 3557 249
rect 3478 173 3557 215
rect 2494 107 2547 173
rect 3500 149 3557 173
rect 3500 115 3512 149
rect 3546 115 3557 149
rect 3500 107 3557 115
rect 3657 249 3714 257
rect 3657 215 3668 249
rect 3702 215 3714 249
rect 3657 149 3714 215
rect 3657 115 3668 149
rect 3702 115 3714 149
rect 3657 107 3714 115
<< mvpdiff >>
rect 801 711 858 719
rect 801 677 813 711
rect 847 677 858 711
rect 801 653 858 677
rect 30 628 83 653
rect 30 594 38 628
rect 72 594 83 628
rect 30 569 83 594
rect 183 628 239 653
rect 183 594 194 628
rect 228 594 239 628
rect 183 569 239 594
rect 339 569 381 653
rect 481 628 537 653
rect 481 594 492 628
rect 526 594 537 628
rect 481 569 537 594
rect 637 569 679 653
rect 779 611 858 653
rect 779 577 813 611
rect 847 577 858 611
rect 779 569 858 577
rect 958 643 1015 719
rect 2178 713 2235 743
rect 958 609 969 643
rect 1003 609 1015 643
rect 958 569 1015 609
rect 1099 675 1156 683
rect 1099 641 1111 675
rect 1145 641 1156 675
rect 1099 575 1156 641
rect 1099 541 1111 575
rect 1145 541 1156 575
rect 1099 533 1156 541
rect 1256 675 1313 683
rect 1256 641 1267 675
rect 1301 641 1313 675
rect 2178 679 2190 713
rect 2224 679 2235 713
rect 1256 575 1313 641
rect 2178 627 2235 679
rect 1256 541 1267 575
rect 1301 541 1313 575
rect 1373 602 1430 627
rect 1373 568 1385 602
rect 1419 568 1430 602
rect 1373 543 1430 568
rect 1530 602 1586 627
rect 1530 568 1541 602
rect 1575 568 1586 602
rect 1530 543 1586 568
rect 1686 543 1728 627
rect 1828 619 1900 627
rect 1828 585 1839 619
rect 1873 585 1900 619
rect 1828 543 1900 585
rect 2000 585 2056 627
rect 2000 551 2011 585
rect 2045 551 2056 585
rect 2000 543 2056 551
rect 2156 543 2235 627
rect 2335 543 2377 743
rect 2477 735 2534 743
rect 2477 701 2488 735
rect 2522 701 2534 735
rect 2477 660 2534 701
rect 2477 626 2488 660
rect 2522 627 2534 660
rect 3067 672 3120 697
rect 3067 638 3075 672
rect 3109 638 3120 672
rect 2522 626 2556 627
rect 2477 585 2556 626
rect 2477 551 2488 585
rect 2522 551 2556 585
rect 2477 543 2556 551
rect 2656 543 2698 627
rect 2798 602 2854 627
rect 2798 568 2809 602
rect 2843 568 2854 602
rect 2798 543 2854 568
rect 2954 602 3007 627
rect 3067 613 3120 638
rect 3220 672 3273 697
rect 3220 638 3231 672
rect 3265 638 3273 672
rect 3508 663 3561 675
rect 3220 613 3273 638
rect 3508 629 3516 663
rect 3550 629 3561 663
rect 3508 625 3561 629
rect 3333 613 3386 625
rect 2954 568 2965 602
rect 2999 568 3007 602
rect 2954 543 3007 568
rect 1256 533 1313 541
rect 3333 579 3341 613
rect 3375 579 3386 613
rect 3333 521 3386 579
rect 3333 487 3341 521
rect 3375 487 3386 521
rect 3333 475 3386 487
rect 3486 592 3561 625
rect 3486 558 3516 592
rect 3550 558 3561 592
rect 3486 521 3561 558
rect 3486 487 3516 521
rect 3550 487 3561 521
rect 3486 475 3561 487
rect 3661 663 3714 675
rect 3661 629 3672 663
rect 3706 629 3714 663
rect 3661 592 3714 629
rect 3661 558 3672 592
rect 3706 558 3714 592
rect 3661 521 3714 558
rect 3661 487 3672 521
rect 3706 487 3714 521
rect 3661 475 3714 487
<< mvndiffc >>
rect 38 132 72 166
rect 194 132 228 166
rect 492 132 526 166
rect 790 132 824 166
rect 946 132 980 166
rect 1056 148 1090 182
rect 1212 148 1246 182
rect 1326 139 1360 173
rect 1482 138 1516 172
rect 1780 138 1814 172
rect 1890 132 1924 166
rect 2207 142 2241 176
rect 2505 195 2539 229
rect 2965 198 2999 232
rect 3154 198 3188 232
rect 3333 198 3367 232
rect 3512 215 3546 249
rect 3512 115 3546 149
rect 3668 215 3702 249
rect 3668 115 3702 149
<< mvpdiffc >>
rect 813 677 847 711
rect 38 594 72 628
rect 194 594 228 628
rect 492 594 526 628
rect 813 577 847 611
rect 969 609 1003 643
rect 1111 641 1145 675
rect 1111 541 1145 575
rect 1267 641 1301 675
rect 2190 679 2224 713
rect 1267 541 1301 575
rect 1385 568 1419 602
rect 1541 568 1575 602
rect 1839 585 1873 619
rect 2011 551 2045 585
rect 2488 701 2522 735
rect 2488 626 2522 660
rect 3075 638 3109 672
rect 2488 551 2522 585
rect 2809 568 2843 602
rect 3231 638 3265 672
rect 3516 629 3550 663
rect 2965 568 2999 602
rect 3341 579 3375 613
rect 3341 487 3375 521
rect 3516 558 3550 592
rect 3516 487 3550 521
rect 3672 629 3706 663
rect 3672 558 3706 592
rect 3672 487 3706 521
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3744 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3744 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 3583 797 3617 831
rect 3679 797 3713 831
<< poly >>
rect 858 719 958 745
rect 2235 743 2335 769
rect 2377 743 2477 769
rect 83 653 183 679
rect 239 653 339 679
rect 381 653 481 679
rect 537 653 637 679
rect 679 653 779 679
rect 1156 683 1256 709
rect 83 547 183 569
rect 239 547 339 569
rect 83 457 339 547
rect 381 471 481 569
rect 537 543 637 569
rect 83 447 239 457
rect 83 417 183 447
rect 83 383 129 417
rect 163 383 183 417
rect 381 437 405 471
rect 439 437 481 471
rect 381 415 481 437
rect 339 403 481 415
rect 339 399 405 403
rect 83 349 183 383
rect 83 315 129 349
rect 163 315 183 349
rect 83 191 183 315
rect 239 369 405 399
rect 439 369 481 403
rect 523 521 637 543
rect 523 487 543 521
rect 577 487 637 521
rect 523 453 637 487
rect 523 419 543 453
rect 577 443 637 453
rect 577 419 623 443
rect 523 399 623 419
rect 239 335 481 369
rect 523 337 637 357
rect 239 191 339 335
rect 523 303 543 337
rect 577 303 637 337
rect 381 263 481 293
rect 381 229 401 263
rect 435 229 481 263
rect 381 191 481 229
rect 523 269 637 303
rect 523 235 543 269
rect 577 235 637 269
rect 523 215 637 235
rect 537 191 637 215
rect 679 353 779 569
rect 858 547 958 569
rect 679 319 700 353
rect 734 319 779 353
rect 679 285 779 319
rect 679 251 700 285
rect 734 251 779 285
rect 679 191 779 251
rect 835 353 958 547
rect 1430 627 1530 653
rect 1586 627 1686 653
rect 1728 627 1828 653
rect 1900 627 2000 653
rect 2056 627 2156 653
rect 3120 697 3220 723
rect 2556 627 2656 653
rect 2698 627 2798 653
rect 2854 627 2954 653
rect 3561 675 3661 701
rect 3386 625 3486 651
rect 1156 511 1256 533
rect 1430 517 1530 543
rect 1586 517 1686 543
rect 835 319 855 353
rect 889 319 958 353
rect 835 285 958 319
rect 835 251 855 285
rect 889 251 958 285
rect 835 217 958 251
rect 1101 477 1256 511
rect 1101 365 1201 477
rect 1298 475 1530 517
rect 1616 495 1686 517
rect 1298 435 1574 475
rect 1616 461 1632 495
rect 1666 461 1686 495
rect 1616 442 1686 461
rect 1728 479 1828 543
rect 1728 445 1774 479
rect 1808 445 1828 479
rect 1101 331 1117 365
rect 1151 331 1201 365
rect 1101 297 1201 331
rect 1101 263 1117 297
rect 1151 263 1201 297
rect 1243 403 1574 435
rect 1243 369 1263 403
rect 1297 400 1574 403
rect 1297 397 1665 400
rect 1297 369 1329 397
rect 1243 335 1329 369
rect 1514 380 1665 397
rect 1243 301 1263 335
rect 1297 301 1329 335
rect 1243 281 1329 301
rect 1371 339 1471 355
rect 1371 305 1412 339
rect 1446 305 1471 339
rect 835 191 935 217
rect 1101 207 1201 263
rect 1371 271 1471 305
rect 1371 237 1412 271
rect 1446 237 1471 271
rect 1371 197 1471 237
rect 1514 346 1611 380
rect 1645 346 1665 380
rect 1514 326 1665 346
rect 1514 223 1627 326
rect 1728 319 1828 445
rect 1900 332 2000 543
rect 2056 521 2156 543
rect 2056 421 2177 521
rect 1728 284 1837 319
rect 1527 197 1627 223
rect 1669 269 1837 284
rect 1669 235 1783 269
rect 1817 235 1837 269
rect 1669 219 1837 235
rect 1900 298 1920 332
rect 1954 313 2000 332
rect 1954 298 2035 313
rect 1669 197 1769 219
rect 1900 213 2035 298
rect 83 81 183 107
rect 239 81 339 107
rect 381 81 481 107
rect 537 81 637 107
rect 679 81 779 107
rect 835 81 935 107
rect 1101 97 1201 123
rect 1935 191 2035 213
rect 2077 269 2177 421
rect 2235 383 2335 543
rect 2377 495 2477 543
rect 2556 521 2656 543
rect 2377 461 2397 495
rect 2431 463 2477 495
rect 2431 461 2451 463
rect 2377 445 2451 461
rect 2519 421 2656 521
rect 2698 521 2798 543
rect 2698 495 2812 521
rect 2698 461 2758 495
rect 2792 461 2812 495
rect 2698 421 2812 461
rect 2493 403 2558 421
rect 2394 387 2558 403
rect 2235 339 2352 383
rect 2235 305 2255 339
rect 2289 305 2352 339
rect 2235 283 2352 305
rect 2077 235 2123 269
rect 2157 235 2177 269
rect 2252 257 2352 283
rect 2394 353 2410 387
rect 2444 362 2558 387
rect 2444 353 2494 362
rect 2394 257 2494 353
rect 2600 333 2670 379
rect 2600 320 2620 333
rect 2569 299 2620 320
rect 2654 299 2670 333
rect 2569 279 2670 299
rect 2569 257 2669 279
rect 2712 257 2812 421
rect 2854 333 2954 543
rect 3120 439 3220 613
rect 2854 299 2870 333
rect 2904 299 2954 333
rect 2854 257 2954 299
rect 3043 419 3220 439
rect 3043 385 3067 419
rect 3101 385 3220 419
rect 3043 383 3220 385
rect 3386 383 3486 475
rect 3561 449 3661 475
rect 3043 351 3486 383
rect 3043 317 3067 351
rect 3101 317 3486 351
rect 3043 283 3486 317
rect 3546 419 3661 449
rect 3546 385 3566 419
rect 3600 385 3661 419
rect 3546 351 3661 385
rect 3546 317 3566 351
rect 3600 317 3661 351
rect 3546 283 3661 317
rect 3043 257 3143 283
rect 3378 257 3478 283
rect 3557 257 3657 283
rect 2077 191 2177 235
rect 1371 87 1471 113
rect 1527 87 1627 113
rect 1669 87 1769 113
rect 2569 147 2669 173
rect 2712 147 2812 173
rect 2854 147 2954 173
rect 3043 147 3143 173
rect 3378 147 3478 173
rect 1935 81 2035 107
rect 2077 81 2177 107
rect 2252 81 2352 107
rect 2394 81 2494 107
rect 3557 81 3657 107
<< polycont >>
rect 129 383 163 417
rect 405 437 439 471
rect 129 315 163 349
rect 405 369 439 403
rect 543 487 577 521
rect 543 419 577 453
rect 543 303 577 337
rect 401 229 435 263
rect 543 235 577 269
rect 700 319 734 353
rect 700 251 734 285
rect 855 319 889 353
rect 855 251 889 285
rect 1632 461 1666 495
rect 1774 445 1808 479
rect 1117 331 1151 365
rect 1117 263 1151 297
rect 1263 369 1297 403
rect 1263 301 1297 335
rect 1412 305 1446 339
rect 1412 237 1446 271
rect 1611 346 1645 380
rect 1783 235 1817 269
rect 1920 298 1954 332
rect 2397 461 2431 495
rect 2758 461 2792 495
rect 2255 305 2289 339
rect 2123 235 2157 269
rect 2410 353 2444 387
rect 2620 299 2654 333
rect 2870 299 2904 333
rect 3067 385 3101 419
rect 3067 317 3101 351
rect 3566 385 3600 419
rect 3566 317 3600 351
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3744 831
rect 124 735 314 741
rect 124 701 130 735
rect 164 701 202 735
rect 236 701 274 735
rect 308 701 314 735
rect 22 628 88 657
rect 22 594 38 628
rect 72 594 88 628
rect 22 541 88 594
rect 124 628 314 701
rect 684 735 863 741
rect 718 701 756 735
rect 790 711 828 735
rect 790 701 813 711
rect 862 701 863 735
rect 684 677 813 701
rect 847 677 863 701
rect 124 594 194 628
rect 228 594 314 628
rect 124 577 314 594
rect 476 628 542 661
rect 476 594 492 628
rect 526 611 542 628
rect 684 611 863 677
rect 526 594 648 611
rect 476 577 648 594
rect 22 521 578 541
rect 22 507 543 521
rect 22 263 56 507
rect 527 487 543 507
rect 577 487 578 521
rect 389 437 405 471
rect 439 437 455 471
rect 113 417 179 433
rect 113 383 129 417
rect 163 383 179 417
rect 113 349 179 383
rect 389 403 455 437
rect 527 453 578 487
rect 527 419 543 453
rect 577 419 578 453
rect 527 403 578 419
rect 614 525 648 577
rect 684 577 813 611
rect 847 577 863 611
rect 684 561 863 577
rect 899 727 1073 761
rect 899 525 933 727
rect 614 491 933 525
rect 969 643 1003 691
rect 389 369 405 403
rect 439 369 455 403
rect 113 315 129 349
rect 163 333 179 349
rect 505 337 578 356
rect 505 333 543 337
rect 163 315 543 333
rect 113 303 543 315
rect 577 303 578 337
rect 113 299 578 303
rect 505 269 578 299
rect 22 229 401 263
rect 435 229 451 263
rect 22 219 451 229
rect 505 235 543 269
rect 577 235 578 269
rect 505 219 578 235
rect 22 166 88 219
rect 614 183 648 491
rect 684 353 750 430
rect 684 319 700 353
rect 734 319 750 353
rect 684 285 750 319
rect 684 251 700 285
rect 734 251 750 285
rect 684 235 750 251
rect 793 353 905 430
rect 793 319 855 353
rect 889 319 905 353
rect 793 285 905 319
rect 793 251 855 285
rect 889 251 905 285
rect 793 235 905 251
rect 969 381 1003 609
rect 1039 489 1073 727
rect 1109 735 1145 741
rect 1109 701 1110 735
rect 1144 701 1145 735
rect 1109 675 1145 701
rect 1109 641 1111 675
rect 1109 575 1145 641
rect 1109 541 1111 575
rect 1109 525 1145 541
rect 1181 727 1419 761
rect 1181 489 1215 727
rect 1039 455 1215 489
rect 1251 675 1306 691
rect 1251 641 1267 675
rect 1301 641 1306 675
rect 1251 575 1306 641
rect 1251 541 1267 575
rect 1301 541 1306 575
rect 1251 419 1306 541
rect 1228 403 1306 419
rect 969 365 1167 381
rect 969 347 1117 365
rect 22 132 38 166
rect 72 132 88 166
rect 22 103 88 132
rect 124 166 314 183
rect 124 132 194 166
rect 228 132 314 166
rect 124 113 314 132
rect 124 79 130 113
rect 164 79 202 113
rect 236 79 274 113
rect 308 79 314 113
rect 476 166 648 183
rect 476 132 492 166
rect 526 149 648 166
rect 684 166 874 199
rect 969 195 1003 347
rect 1101 331 1117 347
rect 1151 331 1167 365
rect 1101 297 1167 331
rect 1101 263 1117 297
rect 1151 263 1167 297
rect 1101 247 1167 263
rect 1228 369 1263 403
rect 1297 369 1306 403
rect 1228 335 1306 369
rect 1228 301 1263 335
rect 1297 301 1306 335
rect 1228 285 1306 301
rect 1342 602 1419 727
rect 1699 735 1889 741
rect 1342 568 1385 602
rect 1342 535 1419 568
rect 1455 671 1661 705
rect 526 132 542 149
rect 476 99 542 132
rect 684 132 790 166
rect 824 132 874 166
rect 684 113 874 132
rect 124 73 314 79
rect 684 79 690 113
rect 724 79 762 113
rect 796 79 834 113
rect 868 79 874 113
rect 930 166 1003 195
rect 930 132 946 166
rect 980 132 1003 166
rect 930 103 1003 132
rect 1040 182 1090 211
rect 1040 148 1056 182
rect 1040 113 1090 148
rect 684 73 874 79
rect 1040 79 1046 113
rect 1080 79 1090 113
rect 1040 73 1090 79
rect 1126 87 1160 247
rect 1228 211 1262 285
rect 1196 182 1262 211
rect 1342 205 1376 535
rect 1455 355 1489 671
rect 1196 148 1212 182
rect 1246 148 1262 182
rect 1196 135 1262 148
rect 1310 173 1376 205
rect 1310 139 1326 173
rect 1360 139 1376 173
rect 1310 123 1376 139
rect 1412 339 1489 355
rect 1446 321 1489 339
rect 1525 602 1591 635
rect 1525 568 1541 602
rect 1575 568 1591 602
rect 1525 535 1591 568
rect 1627 549 1661 671
rect 1699 701 1705 735
rect 1739 701 1777 735
rect 1811 701 1849 735
rect 1883 701 1889 735
rect 1699 619 1889 701
rect 2167 735 2357 751
rect 2167 701 2173 735
rect 2207 713 2245 735
rect 2224 701 2245 713
rect 2279 701 2317 735
rect 2351 701 2357 735
rect 2167 679 2190 701
rect 2224 679 2357 701
rect 2167 657 2357 679
rect 2472 735 2538 751
rect 2472 701 2488 735
rect 2522 701 2538 735
rect 2472 660 2538 701
rect 1699 585 1839 619
rect 1873 585 1889 619
rect 1925 621 2131 655
rect 2472 626 2488 660
rect 2522 626 2538 660
rect 1925 549 1959 621
rect 2097 587 2436 621
rect 1412 271 1446 305
rect 1412 87 1446 237
rect 1525 305 1559 535
rect 1627 515 1959 549
rect 1995 551 2011 585
rect 2045 551 2061 585
rect 1627 495 1682 515
rect 1627 461 1632 495
rect 1666 461 1682 495
rect 1995 479 2061 551
rect 1627 445 1682 461
rect 1758 445 1774 479
rect 1808 445 2061 479
rect 2381 495 2436 587
rect 2472 585 2538 626
rect 2472 551 2488 585
rect 2522 569 2538 585
rect 2653 735 2843 741
rect 2653 701 2659 735
rect 2693 701 2731 735
rect 2765 701 2803 735
rect 2837 701 2843 735
rect 3163 735 3281 741
rect 3163 701 3169 735
rect 3203 701 3241 735
rect 3275 701 3281 735
rect 2653 602 2843 701
rect 2522 551 2584 569
rect 2472 535 2584 551
rect 2653 568 2809 602
rect 2653 535 2843 568
rect 2879 672 3125 701
rect 2879 667 3075 672
rect 2381 461 2397 495
rect 2431 479 2436 495
rect 2431 461 2514 479
rect 2381 445 2514 461
rect 1595 387 2444 409
rect 1595 380 2410 387
rect 1595 346 1611 380
rect 1645 375 2410 380
rect 1645 346 1661 375
rect 1595 341 1661 346
rect 2394 353 2410 375
rect 1697 332 2255 339
rect 1697 305 1920 332
rect 1525 271 1731 305
rect 1904 298 1920 305
rect 1954 305 2255 332
rect 2289 305 2305 339
rect 2394 337 2444 353
rect 1954 298 1970 305
rect 2480 301 2514 445
rect 1904 291 1970 298
rect 1525 205 1559 271
rect 1767 235 1783 269
rect 1817 255 1833 269
rect 1817 235 1940 255
rect 2107 235 2123 269
rect 2157 235 2327 269
rect 1767 221 1940 235
rect 1482 172 1559 205
rect 1516 138 1559 172
rect 1482 105 1559 138
rect 1640 172 1830 185
rect 1640 138 1780 172
rect 1814 138 1830 172
rect 1640 113 1830 138
rect 1126 53 1446 87
rect 1640 79 1646 113
rect 1680 79 1718 113
rect 1752 79 1790 113
rect 1824 79 1830 113
rect 1874 166 1940 221
rect 1874 132 1890 166
rect 1924 132 1940 166
rect 1874 103 1940 132
rect 2067 176 2257 199
rect 2067 142 2207 176
rect 2241 142 2257 176
rect 2067 113 2257 142
rect 1640 73 1830 79
rect 2067 79 2073 113
rect 2107 79 2145 113
rect 2179 79 2217 113
rect 2251 79 2257 113
rect 2067 73 2257 79
rect 2293 87 2327 235
rect 2419 267 2514 301
rect 2550 422 2584 535
rect 2879 499 2913 667
rect 3059 638 3075 667
rect 3109 638 3125 672
rect 2742 495 2913 499
rect 2742 461 2758 495
rect 2792 461 2913 495
rect 2742 458 2913 461
rect 2949 602 3015 631
rect 2949 568 2965 602
rect 2999 568 3015 602
rect 2949 435 3015 568
rect 3059 573 3125 638
rect 3163 672 3281 701
rect 3163 638 3231 672
rect 3265 638 3281 672
rect 3163 609 3281 638
rect 3427 735 3616 741
rect 3427 701 3432 735
rect 3466 701 3504 735
rect 3538 701 3576 735
rect 3610 701 3616 735
rect 3427 663 3616 701
rect 3427 629 3516 663
rect 3550 629 3616 663
rect 3317 613 3391 629
rect 3317 579 3341 613
rect 3375 579 3391 613
rect 3059 539 3204 573
rect 2949 422 3117 435
rect 2550 419 3117 422
rect 2550 388 3067 419
rect 2419 157 2453 267
rect 2550 231 2584 388
rect 3051 385 3067 388
rect 3101 385 3117 419
rect 2489 229 2584 231
rect 2489 195 2505 229
rect 2539 195 2584 229
rect 2489 193 2584 195
rect 2620 333 2670 349
rect 2654 299 2670 333
rect 2620 157 2670 299
rect 2419 123 2670 157
rect 2809 333 2904 352
rect 2809 299 2870 333
rect 3051 351 3117 385
rect 3051 317 3067 351
rect 3101 317 3117 351
rect 3051 301 3117 317
rect 2809 162 2904 299
rect 2940 232 3118 265
rect 2940 198 2965 232
rect 2999 198 3118 232
rect 2809 87 2843 162
rect 2293 53 2843 87
rect 2940 113 3118 198
rect 3154 232 3204 539
rect 3188 198 3204 232
rect 3154 165 3204 198
rect 3317 521 3391 579
rect 3317 487 3341 521
rect 3375 487 3391 521
rect 3317 471 3391 487
rect 3427 592 3616 629
rect 3427 558 3516 592
rect 3550 558 3616 592
rect 3427 521 3616 558
rect 3427 487 3516 521
rect 3550 487 3616 521
rect 3427 471 3616 487
rect 3652 663 3722 679
rect 3652 629 3672 663
rect 3706 629 3722 663
rect 3652 592 3722 629
rect 3652 558 3672 592
rect 3706 558 3722 592
rect 3652 521 3722 558
rect 3652 487 3672 521
rect 3706 487 3722 521
rect 3317 335 3383 471
rect 3550 419 3616 435
rect 3550 385 3566 419
rect 3600 385 3616 419
rect 3550 351 3616 385
rect 3550 335 3566 351
rect 3317 317 3566 335
rect 3600 317 3616 351
rect 3317 301 3616 317
rect 3317 232 3383 301
rect 3317 198 3333 232
rect 3367 198 3383 232
rect 3317 165 3383 198
rect 3419 249 3609 265
rect 3419 215 3512 249
rect 3546 215 3609 249
rect 2974 79 3012 113
rect 3046 79 3084 113
rect 2940 73 3118 79
rect 3419 149 3609 215
rect 3419 115 3512 149
rect 3546 115 3609 149
rect 3419 113 3609 115
rect 3419 79 3425 113
rect 3459 79 3497 113
rect 3531 79 3569 113
rect 3603 79 3609 113
rect 3652 249 3722 487
rect 3652 215 3668 249
rect 3702 215 3722 249
rect 3652 149 3722 215
rect 3652 115 3668 149
rect 3702 115 3722 149
rect 3652 99 3722 115
rect 3419 73 3609 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3744 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 3583 797 3617 831
rect 3679 797 3713 831
rect 130 701 164 735
rect 202 701 236 735
rect 274 701 308 735
rect 684 701 718 735
rect 756 701 790 735
rect 828 711 862 735
rect 828 701 847 711
rect 847 701 862 711
rect 1110 701 1144 735
rect 130 79 164 113
rect 202 79 236 113
rect 274 79 308 113
rect 690 79 724 113
rect 762 79 796 113
rect 834 79 868 113
rect 1046 79 1080 113
rect 1705 701 1739 735
rect 1777 701 1811 735
rect 1849 701 1883 735
rect 2173 713 2207 735
rect 2173 701 2190 713
rect 2190 701 2207 713
rect 2245 701 2279 735
rect 2317 701 2351 735
rect 2659 701 2693 735
rect 2731 701 2765 735
rect 2803 701 2837 735
rect 3169 701 3203 735
rect 3241 701 3275 735
rect 1646 79 1680 113
rect 1718 79 1752 113
rect 1790 79 1824 113
rect 2073 79 2107 113
rect 2145 79 2179 113
rect 2217 79 2251 113
rect 3432 701 3466 735
rect 3504 701 3538 735
rect 3576 701 3610 735
rect 2940 79 2974 113
rect 3012 79 3046 113
rect 3084 79 3118 113
rect 3425 79 3459 113
rect 3497 79 3531 113
rect 3569 79 3603 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
<< metal1 >>
rect 0 831 3744 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3744 831
rect 0 791 3744 797
rect 0 735 3744 763
rect 0 701 130 735
rect 164 701 202 735
rect 236 701 274 735
rect 308 701 684 735
rect 718 701 756 735
rect 790 701 828 735
rect 862 701 1110 735
rect 1144 701 1705 735
rect 1739 701 1777 735
rect 1811 701 1849 735
rect 1883 701 2173 735
rect 2207 701 2245 735
rect 2279 701 2317 735
rect 2351 701 2659 735
rect 2693 701 2731 735
rect 2765 701 2803 735
rect 2837 701 3169 735
rect 3203 701 3241 735
rect 3275 701 3432 735
rect 3466 701 3504 735
rect 3538 701 3576 735
rect 3610 701 3744 735
rect 0 689 3744 701
rect 0 113 3744 125
rect 0 79 130 113
rect 164 79 202 113
rect 236 79 274 113
rect 308 79 690 113
rect 724 79 762 113
rect 796 79 834 113
rect 868 79 1046 113
rect 1080 79 1646 113
rect 1680 79 1718 113
rect 1752 79 1790 113
rect 1824 79 2073 113
rect 2107 79 2145 113
rect 2179 79 2217 113
rect 2251 79 2940 113
rect 2974 79 3012 113
rect 3046 79 3084 113
rect 3118 79 3425 113
rect 3459 79 3497 113
rect 3531 79 3569 113
rect 3603 79 3744 113
rect 0 51 3744 79
rect 0 17 3744 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3744 17
rect 0 -23 3744 -17
<< labels >>
flabel comment s 1776 362 1776 362 0 FreeSans 200 90 0 0 no_jumper_check
flabel comment s 1435 420 1435 420 0 FreeSans 200 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 sdfstp_1
flabel metal1 s 0 51 3744 125 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel metal1 s 0 0 3744 23 0 FreeSans 340 0 0 0 VNB
port 7 nsew ground bidirectional
flabel metal1 s 0 689 3744 763 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 791 3744 814 0 FreeSans 340 0 0 0 VPB
port 8 nsew power bidirectional
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 3679 168 3713 202 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3679 242 3713 276 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3679 316 3713 350 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3679 390 3713 424 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3679 464 3713 498 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3679 538 3713 572 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3679 612 3713 646 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2815 168 2849 202 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 2815 242 2849 276 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 2815 316 2849 350 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
rlabel locali s 2067 73 2257 199 1 VGND
port 6 nsew ground bidirectional
rlabel locali s 2940 73 3118 265 1 VGND
port 6 nsew ground bidirectional
rlabel locali s 3419 73 3609 265 1 VGND
port 6 nsew ground bidirectional
rlabel locali s 684 73 874 199 1 VGND
port 6 nsew ground bidirectional
rlabel locali s 1040 73 1090 211 1 VGND
port 6 nsew ground bidirectional
rlabel locali s 1640 73 1830 185 1 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 51 3744 125 1 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 -23 3744 23 1 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 791 3744 837 1 VPB
port 8 nsew power bidirectional
rlabel locali s 2167 657 2357 751 1 VPWR
port 9 nsew power bidirectional
rlabel locali s 2653 535 2843 741 1 VPWR
port 9 nsew power bidirectional
rlabel locali s 3163 609 3281 741 1 VPWR
port 9 nsew power bidirectional
rlabel locali s 3427 471 3616 741 1 VPWR
port 9 nsew power bidirectional
rlabel locali s 684 561 863 741 1 VPWR
port 9 nsew power bidirectional
rlabel locali s 1109 525 1145 741 1 VPWR
port 9 nsew power bidirectional
rlabel locali s 1699 585 1889 741 1 VPWR
port 9 nsew power bidirectional
rlabel metal1 s 0 689 3744 763 1 VPWR
port 9 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 3744 814
string GDS_END 605350
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 570398
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
