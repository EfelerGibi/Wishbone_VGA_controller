magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 99 157 509 203
rect 1 21 721 157
rect 29 -17 63 21
<< locali >>
rect 17 199 99 323
rect 554 325 619 492
rect 573 255 619 325
rect 573 153 719 255
rect 573 123 619 153
rect 554 57 619 123
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 19 391 69 493
rect 115 425 181 527
rect 19 357 167 391
rect 133 350 167 357
rect 133 265 201 350
rect 235 285 288 493
rect 339 349 389 493
rect 427 383 493 527
rect 339 300 519 349
rect 653 327 719 527
rect 241 265 288 285
rect 133 199 207 265
rect 241 199 433 265
rect 133 162 168 199
rect 19 128 168 162
rect 241 156 285 199
rect 467 161 519 300
rect 19 61 69 128
rect 115 17 181 94
rect 219 51 285 156
rect 323 127 519 161
rect 323 51 389 127
rect 427 17 493 93
rect 653 17 719 110
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 17 199 99 323 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 736 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 1 21 721 157 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 99 157 509 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 554 57 619 123 6 X
port 6 nsew signal output
rlabel locali s 573 123 619 153 6 X
port 6 nsew signal output
rlabel locali s 573 153 719 255 6 X
port 6 nsew signal output
rlabel locali s 573 255 619 325 6 X
port 6 nsew signal output
rlabel locali s 554 325 619 492 6 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 736 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3290926
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3284314
<< end >>
