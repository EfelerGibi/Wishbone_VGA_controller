magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect 0 0 642 708
<< pmos >>
rect 171 189 201 519
rect 257 189 293 519
rect 349 189 385 519
rect 441 189 471 519
<< pdiff >>
rect 111 507 171 519
rect 111 473 126 507
rect 160 473 171 507
rect 111 439 171 473
rect 111 405 126 439
rect 160 405 171 439
rect 111 371 171 405
rect 111 337 126 371
rect 160 337 171 371
rect 111 303 171 337
rect 111 269 126 303
rect 160 269 171 303
rect 111 235 171 269
rect 111 201 126 235
rect 160 201 171 235
rect 111 189 171 201
rect 201 507 257 519
rect 201 473 212 507
rect 246 473 257 507
rect 201 439 257 473
rect 201 405 212 439
rect 246 405 257 439
rect 201 371 257 405
rect 201 337 212 371
rect 246 337 257 371
rect 201 303 257 337
rect 201 269 212 303
rect 246 269 257 303
rect 201 235 257 269
rect 201 201 212 235
rect 246 201 257 235
rect 201 189 257 201
rect 293 507 349 519
rect 293 473 304 507
rect 338 473 349 507
rect 293 439 349 473
rect 293 405 304 439
rect 338 405 349 439
rect 293 371 349 405
rect 293 337 304 371
rect 338 337 349 371
rect 293 303 349 337
rect 293 269 304 303
rect 338 269 349 303
rect 293 235 349 269
rect 293 201 304 235
rect 338 201 349 235
rect 293 189 349 201
rect 385 507 441 519
rect 385 473 396 507
rect 430 473 441 507
rect 385 439 441 473
rect 385 405 396 439
rect 430 405 441 439
rect 385 371 441 405
rect 385 337 396 371
rect 430 337 441 371
rect 385 303 441 337
rect 385 269 396 303
rect 430 269 441 303
rect 385 235 441 269
rect 385 201 396 235
rect 430 201 441 235
rect 385 189 441 201
rect 471 507 531 519
rect 471 473 482 507
rect 516 473 531 507
rect 471 439 531 473
rect 471 405 482 439
rect 516 405 531 439
rect 471 371 531 405
rect 471 337 482 371
rect 516 337 531 371
rect 471 303 531 337
rect 471 269 482 303
rect 516 269 531 303
rect 471 235 531 269
rect 471 201 482 235
rect 516 201 531 235
rect 471 189 531 201
<< pdiffc >>
rect 126 473 160 507
rect 126 405 160 439
rect 126 337 160 371
rect 126 269 160 303
rect 126 201 160 235
rect 212 473 246 507
rect 212 405 246 439
rect 212 337 246 371
rect 212 269 246 303
rect 212 201 246 235
rect 304 473 338 507
rect 304 405 338 439
rect 304 337 338 371
rect 304 269 338 303
rect 304 201 338 235
rect 396 473 430 507
rect 396 405 430 439
rect 396 337 430 371
rect 396 269 430 303
rect 396 201 430 235
rect 482 473 516 507
rect 482 405 516 439
rect 482 337 516 371
rect 482 269 516 303
rect 482 201 516 235
<< nsubdiff >>
rect 41 507 111 519
rect 41 473 58 507
rect 92 473 111 507
rect 41 439 111 473
rect 41 405 58 439
rect 92 405 111 439
rect 41 371 111 405
rect 41 337 58 371
rect 92 337 111 371
rect 41 303 111 337
rect 41 269 58 303
rect 92 269 111 303
rect 41 235 111 269
rect 41 201 58 235
rect 92 201 111 235
rect 41 189 111 201
rect 531 507 601 519
rect 531 473 550 507
rect 584 473 601 507
rect 531 439 601 473
rect 531 405 550 439
rect 584 405 601 439
rect 531 371 601 405
rect 531 337 550 371
rect 584 337 601 371
rect 531 303 601 337
rect 531 269 550 303
rect 584 269 601 303
rect 531 235 601 269
rect 531 201 550 235
rect 584 201 601 235
rect 531 189 601 201
<< nsubdiffcont >>
rect 58 473 92 507
rect 58 405 92 439
rect 58 337 92 371
rect 58 269 92 303
rect 58 201 92 235
rect 550 473 584 507
rect 550 405 584 439
rect 550 337 584 371
rect 550 269 584 303
rect 550 201 584 235
<< poly >>
rect 243 687 399 708
rect 243 653 264 687
rect 298 653 344 687
rect 378 653 399 687
rect 243 619 399 653
rect 120 601 201 617
rect 120 567 136 601
rect 170 567 201 601
rect 243 585 264 619
rect 298 585 344 619
rect 378 585 399 619
rect 243 569 399 585
rect 441 601 522 617
rect 120 551 201 567
rect 171 519 201 551
rect 257 519 293 569
rect 349 519 385 569
rect 441 567 472 601
rect 506 567 522 601
rect 441 551 522 567
rect 441 519 471 551
rect 171 157 201 189
rect 120 141 201 157
rect 120 107 136 141
rect 170 107 201 141
rect 257 139 293 189
rect 349 139 385 189
rect 441 157 471 189
rect 441 141 522 157
rect 120 91 201 107
rect 243 123 399 139
rect 243 89 264 123
rect 298 89 344 123
rect 378 89 399 123
rect 441 107 472 141
rect 506 107 522 141
rect 441 91 522 107
rect 243 55 399 89
rect 243 21 264 55
rect 298 21 344 55
rect 378 21 399 55
rect 243 0 399 21
<< polycont >>
rect 264 653 298 687
rect 344 653 378 687
rect 136 567 170 601
rect 264 585 298 619
rect 344 585 378 619
rect 472 567 506 601
rect 136 107 170 141
rect 264 89 298 123
rect 344 89 378 123
rect 472 107 506 141
rect 264 21 298 55
rect 344 21 378 55
<< locali >>
rect 248 689 394 708
rect 248 655 262 689
rect 296 687 346 689
rect 248 653 264 655
rect 298 653 344 687
rect 380 655 394 689
rect 378 653 394 655
rect 248 619 394 653
rect 248 617 264 619
rect 120 601 186 617
rect 120 567 136 601
rect 170 567 186 601
rect 248 583 262 617
rect 298 585 344 619
rect 378 617 394 619
rect 296 583 346 585
rect 380 583 394 617
rect 248 569 394 583
rect 456 601 522 617
rect 120 551 186 567
rect 456 567 472 601
rect 506 567 522 601
rect 456 551 522 567
rect 120 523 160 551
rect 482 523 522 551
rect 41 507 160 523
rect 41 473 58 507
rect 92 479 126 507
rect 94 473 126 479
rect 41 445 60 473
rect 94 445 160 473
rect 41 439 160 445
rect 41 405 58 439
rect 92 407 126 439
rect 94 405 126 407
rect 41 373 60 405
rect 94 373 160 405
rect 41 371 160 373
rect 41 337 58 371
rect 92 337 126 371
rect 41 335 160 337
rect 41 303 60 335
rect 94 303 160 335
rect 41 269 58 303
rect 94 301 126 303
rect 92 269 126 301
rect 41 263 160 269
rect 41 235 60 263
rect 94 235 160 263
rect 41 201 58 235
rect 94 229 126 235
rect 92 201 126 229
rect 41 185 160 201
rect 212 507 246 523
rect 212 439 246 445
rect 212 371 246 373
rect 212 335 246 337
rect 212 263 246 269
rect 212 185 246 201
rect 304 507 338 523
rect 304 439 338 445
rect 304 371 338 373
rect 304 335 338 337
rect 304 263 338 269
rect 304 185 338 201
rect 396 507 430 523
rect 396 439 430 445
rect 396 371 430 373
rect 396 335 430 337
rect 396 263 430 269
rect 396 185 430 201
rect 482 507 601 523
rect 516 479 550 507
rect 516 473 548 479
rect 584 473 601 507
rect 482 445 548 473
rect 582 445 601 473
rect 482 439 601 445
rect 516 407 550 439
rect 516 405 548 407
rect 584 405 601 439
rect 482 373 548 405
rect 582 373 601 405
rect 482 371 601 373
rect 516 337 550 371
rect 584 337 601 371
rect 482 335 601 337
rect 482 303 548 335
rect 582 303 601 335
rect 516 301 548 303
rect 516 269 550 301
rect 584 269 601 303
rect 482 263 601 269
rect 482 235 548 263
rect 582 235 601 263
rect 516 229 548 235
rect 516 201 550 229
rect 584 201 601 235
rect 482 185 601 201
rect 120 157 160 185
rect 482 157 522 185
rect 120 141 186 157
rect 120 107 136 141
rect 170 107 186 141
rect 456 141 522 157
rect 120 91 186 107
rect 248 125 394 139
rect 248 91 262 125
rect 296 123 346 125
rect 248 89 264 91
rect 298 89 344 123
rect 380 91 394 125
rect 456 107 472 141
rect 506 107 522 141
rect 456 91 522 107
rect 378 89 394 91
rect 248 55 394 89
rect 248 53 264 55
rect 248 19 262 53
rect 298 21 344 55
rect 378 53 394 55
rect 296 19 346 21
rect 380 19 394 53
rect 248 0 394 19
<< viali >>
rect 262 687 296 689
rect 346 687 380 689
rect 262 655 264 687
rect 264 655 296 687
rect 346 655 378 687
rect 378 655 380 687
rect 262 585 264 617
rect 264 585 296 617
rect 346 585 378 617
rect 378 585 380 617
rect 262 583 296 585
rect 346 583 380 585
rect 60 473 92 479
rect 92 473 94 479
rect 60 445 94 473
rect 60 405 92 407
rect 92 405 94 407
rect 60 373 94 405
rect 60 303 94 335
rect 60 301 92 303
rect 92 301 94 303
rect 60 235 94 263
rect 60 229 92 235
rect 92 229 94 235
rect 212 473 246 479
rect 212 445 246 473
rect 212 405 246 407
rect 212 373 246 405
rect 212 303 246 335
rect 212 301 246 303
rect 212 235 246 263
rect 212 229 246 235
rect 304 473 338 479
rect 304 445 338 473
rect 304 405 338 407
rect 304 373 338 405
rect 304 303 338 335
rect 304 301 338 303
rect 304 235 338 263
rect 304 229 338 235
rect 396 473 430 479
rect 396 445 430 473
rect 396 405 430 407
rect 396 373 430 405
rect 396 303 430 335
rect 396 301 430 303
rect 396 235 430 263
rect 396 229 430 235
rect 548 473 550 479
rect 550 473 582 479
rect 548 445 582 473
rect 548 405 550 407
rect 550 405 582 407
rect 548 373 582 405
rect 548 303 582 335
rect 548 301 550 303
rect 550 301 582 303
rect 548 235 582 263
rect 548 229 550 235
rect 550 229 582 235
rect 262 123 296 125
rect 346 123 380 125
rect 262 91 264 123
rect 264 91 296 123
rect 346 91 378 123
rect 378 91 380 123
rect 262 21 264 53
rect 264 21 296 53
rect 346 21 378 53
rect 378 21 380 53
rect 262 19 296 21
rect 346 19 380 21
<< metal1 >>
rect 250 689 392 708
rect 250 655 262 689
rect 296 655 346 689
rect 380 655 392 689
rect 250 617 392 655
rect 250 583 262 617
rect 296 583 346 617
rect 380 583 392 617
rect 250 571 392 583
rect 41 479 100 507
rect 41 445 60 479
rect 94 445 100 479
rect 41 407 100 445
rect 41 373 60 407
rect 94 373 100 407
rect 41 335 100 373
rect 41 301 60 335
rect 94 301 100 335
rect 41 263 100 301
rect 41 229 60 263
rect 94 229 100 263
rect 41 201 100 229
rect 203 479 255 507
rect 203 445 212 479
rect 246 445 255 479
rect 203 407 255 445
rect 203 373 212 407
rect 246 373 255 407
rect 203 335 255 373
rect 203 323 212 335
rect 246 323 255 335
rect 203 263 255 271
rect 203 259 212 263
rect 246 259 255 263
rect 203 201 255 207
rect 295 501 347 507
rect 295 445 304 449
rect 338 445 347 449
rect 295 437 347 445
rect 295 373 304 385
rect 338 373 347 385
rect 295 335 347 373
rect 295 301 304 335
rect 338 301 347 335
rect 295 263 347 301
rect 295 229 304 263
rect 338 229 347 263
rect 295 201 347 229
rect 387 479 439 507
rect 387 445 396 479
rect 430 445 439 479
rect 387 407 439 445
rect 387 373 396 407
rect 430 373 439 407
rect 387 335 439 373
rect 387 323 396 335
rect 430 323 439 335
rect 387 263 439 271
rect 387 259 396 263
rect 430 259 439 263
rect 387 201 439 207
rect 542 479 601 507
rect 542 445 548 479
rect 582 445 601 479
rect 542 407 601 445
rect 542 373 548 407
rect 582 373 601 407
rect 542 335 601 373
rect 542 301 548 335
rect 582 301 601 335
rect 542 263 601 301
rect 542 229 548 263
rect 582 229 601 263
rect 542 201 601 229
rect 250 125 392 137
rect 250 91 262 125
rect 296 91 346 125
rect 380 91 392 125
rect 250 53 392 91
rect 250 19 262 53
rect 296 19 346 53
rect 380 19 392 53
rect 250 0 392 19
<< via1 >>
rect 203 301 212 323
rect 212 301 246 323
rect 246 301 255 323
rect 203 271 255 301
rect 203 229 212 259
rect 212 229 246 259
rect 246 229 255 259
rect 203 207 255 229
rect 295 479 347 501
rect 295 449 304 479
rect 304 449 338 479
rect 338 449 347 479
rect 295 407 347 437
rect 295 385 304 407
rect 304 385 338 407
rect 338 385 347 407
rect 387 301 396 323
rect 396 301 430 323
rect 430 301 439 323
rect 387 271 439 301
rect 387 229 396 259
rect 396 229 430 259
rect 430 229 439 259
rect 387 207 439 229
<< metal2 >>
rect 14 501 628 507
rect 14 449 295 501
rect 347 449 628 501
rect 14 437 628 449
rect 14 385 295 437
rect 347 385 628 437
rect 14 379 628 385
rect 14 323 628 329
rect 14 271 203 323
rect 255 271 387 323
rect 439 271 628 323
rect 14 259 628 271
rect 14 207 203 259
rect 255 207 387 259
rect 439 207 628 259
rect 14 201 628 207
<< labels >>
flabel comment s 184 343 184 343 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 453 344 453 344 0 FreeSans 180 90 0 0 dummy_poly
flabel metal1 s 255 608 386 659 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal1 s 255 44 386 95 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal1 s 41 339 87 369 0 FreeSans 200 90 0 0 BULK
port 4 nsew
flabel metal1 s 555 339 601 369 0 FreeSans 200 90 0 0 BULK
port 4 nsew
flabel metal2 s 14 201 35 329 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal2 s 14 379 35 507 7 FreeSans 300 180 0 0 DRAIN
port 1 nsew
<< properties >>
string GDS_END 9474790
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9463698
string device primitive
<< end >>
