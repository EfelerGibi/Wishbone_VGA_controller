magic
tech sky130A
magscale 1 2
timestamp 1685806364
<< nwell >>
rect 1066 349509 558846 349830
rect 1066 348421 558846 348987
rect 1066 347333 558846 347899
rect 1066 346245 558846 346811
rect 1066 345157 558846 345723
rect 1066 344069 558846 344635
rect 1066 342981 558846 343547
rect 1066 341893 558846 342459
rect 1066 340805 558846 341371
rect 1066 339717 558846 340283
rect 1066 338629 558846 339195
rect 1066 337541 558846 338107
rect 1066 336453 558846 337019
rect 1066 335365 558846 335931
rect 1066 334277 558846 334843
rect 1066 333189 558846 333755
rect 1066 332101 558846 332667
rect 1066 331013 558846 331579
rect 1066 329925 558846 330491
rect 1066 328837 558846 329403
rect 1066 327749 558846 328315
rect 1066 326661 558846 327227
rect 1066 325573 558846 326139
rect 1066 324485 558846 325051
rect 1066 323397 558846 323963
rect 1066 322309 558846 322875
rect 1066 321221 558846 321787
rect 1066 320133 558846 320699
rect 1066 319045 558846 319611
rect 1066 317957 558846 318523
rect 1066 316869 558846 317435
rect 1066 315781 558846 316347
rect 1066 314693 558846 315259
rect 1066 313605 558846 314171
rect 1066 312517 558846 313083
rect 1066 311429 558846 311995
rect 1066 310341 558846 310907
rect 1066 309253 558846 309819
rect 1066 308165 558846 308731
rect 1066 307077 558846 307643
rect 1066 305989 558846 306555
rect 1066 304901 558846 305467
rect 1066 303813 558846 304379
rect 1066 302725 558846 303291
rect 1066 301637 558846 302203
rect 1066 300549 558846 301115
rect 1066 299461 558846 300027
rect 1066 298373 558846 298939
rect 1066 297285 558846 297851
rect 1066 296197 558846 296763
rect 1066 295109 558846 295675
rect 1066 294021 558846 294587
rect 1066 292933 558846 293499
rect 1066 291845 558846 292411
rect 1066 290757 558846 291323
rect 1066 289669 558846 290235
rect 1066 288581 558846 289147
rect 1066 287493 558846 288059
rect 1066 286405 558846 286971
rect 1066 285317 558846 285883
rect 1066 284229 558846 284795
rect 1066 283141 558846 283707
rect 1066 282053 558846 282619
rect 1066 280965 558846 281531
rect 1066 279877 558846 280443
rect 1066 278789 558846 279355
rect 1066 277701 558846 278267
rect 1066 276613 558846 277179
rect 1066 275525 558846 276091
rect 1066 274437 558846 275003
rect 1066 273349 558846 273915
rect 1066 272261 558846 272827
rect 1066 271173 558846 271739
rect 1066 270085 558846 270651
rect 1066 268997 558846 269563
rect 1066 267909 558846 268475
rect 1066 266821 558846 267387
rect 1066 265733 558846 266299
rect 1066 264645 558846 265211
rect 1066 263557 558846 264123
rect 1066 262469 558846 263035
rect 1066 261381 558846 261947
rect 1066 260293 558846 260859
rect 1066 259205 558846 259771
rect 1066 258117 558846 258683
rect 1066 257029 558846 257595
rect 1066 255941 558846 256507
rect 1066 254853 558846 255419
rect 1066 253765 558846 254331
rect 1066 252677 558846 253243
rect 1066 251589 558846 252155
rect 1066 250501 558846 251067
rect 1066 249413 558846 249979
rect 1066 248325 558846 248891
rect 1066 247237 558846 247803
rect 1066 246149 558846 246715
rect 1066 245061 558846 245627
rect 1066 243973 558846 244539
rect 1066 242885 558846 243451
rect 1066 241797 558846 242363
rect 1066 240709 558846 241275
rect 1066 239621 558846 240187
rect 1066 238533 558846 239099
rect 1066 237445 558846 238011
rect 1066 236357 558846 236923
rect 1066 235269 558846 235835
rect 1066 234181 558846 234747
rect 1066 233093 558846 233659
rect 1066 232005 558846 232571
rect 1066 230917 558846 231483
rect 1066 229829 558846 230395
rect 1066 228741 558846 229307
rect 1066 227653 558846 228219
rect 1066 226565 558846 227131
rect 1066 225477 558846 226043
rect 1066 224389 558846 224955
rect 1066 223301 558846 223867
rect 1066 222213 558846 222779
rect 1066 221125 558846 221691
rect 1066 220037 558846 220603
rect 1066 218949 558846 219515
rect 1066 217861 558846 218427
rect 1066 216773 558846 217339
rect 1066 215685 558846 216251
rect 1066 214597 558846 215163
rect 1066 213509 558846 214075
rect 1066 212421 558846 212987
rect 1066 211333 558846 211899
rect 1066 210245 558846 210811
rect 1066 209157 558846 209723
rect 1066 208069 558846 208635
rect 1066 206981 558846 207547
rect 1066 205893 558846 206459
rect 1066 204805 558846 205371
rect 1066 203717 558846 204283
rect 1066 202629 558846 203195
rect 1066 201541 558846 202107
rect 1066 200453 558846 201019
rect 1066 199365 558846 199931
rect 1066 198277 558846 198843
rect 1066 197189 558846 197755
rect 1066 196101 558846 196667
rect 1066 195013 558846 195579
rect 1066 193925 558846 194491
rect 1066 192837 558846 193403
rect 1066 191749 558846 192315
rect 1066 190661 558846 191227
rect 1066 189573 558846 190139
rect 1066 188485 558846 189051
rect 1066 187397 558846 187963
rect 1066 186309 558846 186875
rect 1066 185221 558846 185787
rect 1066 184133 558846 184699
rect 1066 183045 558846 183611
rect 1066 181957 558846 182523
rect 1066 180869 558846 181435
rect 1066 179781 558846 180347
rect 1066 178693 558846 179259
rect 1066 177605 558846 178171
rect 1066 176517 558846 177083
rect 1066 175429 558846 175995
rect 1066 174341 558846 174907
rect 1066 173253 558846 173819
rect 1066 172165 558846 172731
rect 1066 171077 558846 171643
rect 1066 169989 558846 170555
rect 1066 168901 558846 169467
rect 1066 167813 558846 168379
rect 1066 166725 558846 167291
rect 1066 165637 558846 166203
rect 1066 164549 558846 165115
rect 1066 163461 558846 164027
rect 1066 162373 558846 162939
rect 1066 161285 558846 161851
rect 1066 160197 558846 160763
rect 1066 159109 558846 159675
rect 1066 158021 558846 158587
rect 1066 156933 558846 157499
rect 1066 155845 558846 156411
rect 1066 154757 558846 155323
rect 1066 153669 558846 154235
rect 1066 152581 558846 153147
rect 1066 151493 558846 152059
rect 1066 150405 558846 150971
rect 1066 149317 558846 149883
rect 1066 148229 558846 148795
rect 1066 147141 558846 147707
rect 1066 146053 558846 146619
rect 1066 144965 558846 145531
rect 1066 143877 558846 144443
rect 1066 142789 558846 143355
rect 1066 141701 558846 142267
rect 1066 140613 558846 141179
rect 1066 139525 558846 140091
rect 1066 138437 558846 139003
rect 1066 137349 558846 137915
rect 1066 136261 558846 136827
rect 1066 135173 558846 135739
rect 1066 134085 558846 134651
rect 1066 132997 558846 133563
rect 1066 131909 558846 132475
rect 1066 130821 558846 131387
rect 1066 129733 558846 130299
rect 1066 128645 558846 129211
rect 1066 127557 558846 128123
rect 1066 126469 558846 127035
rect 1066 125381 558846 125947
rect 1066 124293 558846 124859
rect 1066 123205 558846 123771
rect 1066 122117 558846 122683
rect 1066 121029 558846 121595
rect 1066 119941 558846 120507
rect 1066 118853 558846 119419
rect 1066 117765 558846 118331
rect 1066 116677 558846 117243
rect 1066 115589 558846 116155
rect 1066 114501 558846 115067
rect 1066 113413 558846 113979
rect 1066 112325 558846 112891
rect 1066 111237 558846 111803
rect 1066 110149 558846 110715
rect 1066 109061 558846 109627
rect 1066 107973 558846 108539
rect 1066 106885 558846 107451
rect 1066 105797 558846 106363
rect 1066 104709 558846 105275
rect 1066 103621 558846 104187
rect 1066 102533 558846 103099
rect 1066 101445 558846 102011
rect 1066 100357 558846 100923
rect 1066 99269 558846 99835
rect 1066 98181 558846 98747
rect 1066 97093 558846 97659
rect 1066 96005 558846 96571
rect 1066 94917 558846 95483
rect 1066 93829 558846 94395
rect 1066 92741 558846 93307
rect 1066 91653 558846 92219
rect 1066 90565 558846 91131
rect 1066 89477 558846 90043
rect 1066 88389 558846 88955
rect 1066 87301 558846 87867
rect 1066 86213 558846 86779
rect 1066 85125 558846 85691
rect 1066 84037 558846 84603
rect 1066 82949 558846 83515
rect 1066 81861 558846 82427
rect 1066 80773 558846 81339
rect 1066 79685 558846 80251
rect 1066 78597 558846 79163
rect 1066 77509 558846 78075
rect 1066 76421 558846 76987
rect 1066 75333 558846 75899
rect 1066 74245 558846 74811
rect 1066 73157 558846 73723
rect 1066 72069 558846 72635
rect 1066 70981 558846 71547
rect 1066 69893 558846 70459
rect 1066 68805 558846 69371
rect 1066 67717 558846 68283
rect 1066 66629 558846 67195
rect 1066 65541 558846 66107
rect 1066 64453 558846 65019
rect 1066 63365 558846 63931
rect 1066 62277 558846 62843
rect 1066 61189 558846 61755
rect 1066 60101 558846 60667
rect 1066 59013 558846 59579
rect 1066 57925 558846 58491
rect 1066 56837 558846 57403
rect 1066 55749 558846 56315
rect 1066 54661 558846 55227
rect 1066 53573 558846 54139
rect 1066 52485 558846 53051
rect 1066 51397 558846 51963
rect 1066 50309 558846 50875
rect 1066 49221 558846 49787
rect 1066 48133 558846 48699
rect 1066 47045 558846 47611
rect 1066 45957 558846 46523
rect 1066 44869 558846 45435
rect 1066 43781 558846 44347
rect 1066 42693 558846 43259
rect 1066 41605 558846 42171
rect 1066 40517 558846 41083
rect 1066 39429 558846 39995
rect 1066 38341 558846 38907
rect 1066 37253 558846 37819
rect 1066 36165 558846 36731
rect 1066 35077 558846 35643
rect 1066 33989 558846 34555
rect 1066 32901 558846 33467
rect 1066 31813 558846 32379
rect 1066 30725 558846 31291
rect 1066 29637 558846 30203
rect 1066 28549 558846 29115
rect 1066 27461 558846 28027
rect 1066 26373 558846 26939
rect 1066 25285 558846 25851
rect 1066 24197 558846 24763
rect 1066 23109 558846 23675
rect 1066 22021 558846 22587
rect 1066 20933 558846 21499
rect 1066 19845 558846 20411
rect 1066 18757 558846 19323
rect 1066 17669 558846 18235
rect 1066 16581 558846 17147
rect 1066 15493 558846 16059
rect 1066 14405 558846 14971
rect 1066 13317 558846 13883
rect 1066 12229 558846 12795
rect 1066 11141 558846 11707
rect 1066 10053 558846 10619
rect 1066 8965 558846 9531
rect 1066 7877 558846 8443
rect 1066 6789 558846 7355
rect 1066 5701 558846 6267
rect 1066 4613 558846 5179
rect 1066 3525 558846 4091
rect 1066 2437 558846 3003
<< obsli1 >>
rect 1104 2159 558808 349809
<< obsm1 >>
rect 1104 552 558808 349840
<< metal2 >>
rect 4894 0 4950 800
rect 9126 0 9182 800
rect 13358 0 13414 800
rect 17590 0 17646 800
rect 21822 0 21878 800
rect 26054 0 26110 800
rect 30286 0 30342 800
rect 34518 0 34574 800
rect 38750 0 38806 800
rect 42982 0 43038 800
rect 47214 0 47270 800
rect 51446 0 51502 800
rect 55678 0 55734 800
rect 59910 0 59966 800
rect 64142 0 64198 800
rect 68374 0 68430 800
rect 72606 0 72662 800
rect 76838 0 76894 800
rect 81070 0 81126 800
rect 85302 0 85358 800
rect 89534 0 89590 800
rect 93766 0 93822 800
rect 97998 0 98054 800
rect 102230 0 102286 800
rect 106462 0 106518 800
rect 110694 0 110750 800
rect 114926 0 114982 800
rect 119158 0 119214 800
rect 123390 0 123446 800
rect 127622 0 127678 800
rect 131854 0 131910 800
rect 136086 0 136142 800
rect 140318 0 140374 800
rect 144550 0 144606 800
rect 148782 0 148838 800
rect 153014 0 153070 800
rect 157246 0 157302 800
rect 161478 0 161534 800
rect 165710 0 165766 800
rect 169942 0 169998 800
rect 174174 0 174230 800
rect 178406 0 178462 800
rect 182638 0 182694 800
rect 186870 0 186926 800
rect 191102 0 191158 800
rect 195334 0 195390 800
rect 199566 0 199622 800
rect 203798 0 203854 800
rect 208030 0 208086 800
rect 212262 0 212318 800
rect 216494 0 216550 800
rect 220726 0 220782 800
rect 224958 0 225014 800
rect 229190 0 229246 800
rect 233422 0 233478 800
rect 237654 0 237710 800
rect 241886 0 241942 800
rect 246118 0 246174 800
rect 250350 0 250406 800
rect 254582 0 254638 800
rect 258814 0 258870 800
rect 263046 0 263102 800
rect 267278 0 267334 800
rect 271510 0 271566 800
rect 275742 0 275798 800
rect 279974 0 280030 800
rect 284206 0 284262 800
rect 288438 0 288494 800
rect 292670 0 292726 800
rect 296902 0 296958 800
rect 301134 0 301190 800
rect 305366 0 305422 800
rect 309598 0 309654 800
rect 313830 0 313886 800
rect 318062 0 318118 800
rect 322294 0 322350 800
rect 326526 0 326582 800
rect 330758 0 330814 800
rect 334990 0 335046 800
rect 339222 0 339278 800
rect 343454 0 343510 800
rect 347686 0 347742 800
rect 351918 0 351974 800
rect 356150 0 356206 800
rect 360382 0 360438 800
rect 364614 0 364670 800
rect 368846 0 368902 800
rect 373078 0 373134 800
rect 377310 0 377366 800
rect 381542 0 381598 800
rect 385774 0 385830 800
rect 390006 0 390062 800
rect 394238 0 394294 800
rect 398470 0 398526 800
rect 402702 0 402758 800
rect 406934 0 406990 800
rect 411166 0 411222 800
rect 415398 0 415454 800
rect 419630 0 419686 800
rect 423862 0 423918 800
rect 428094 0 428150 800
rect 432326 0 432382 800
rect 436558 0 436614 800
rect 440790 0 440846 800
rect 445022 0 445078 800
rect 449254 0 449310 800
rect 453486 0 453542 800
rect 457718 0 457774 800
rect 461950 0 462006 800
rect 466182 0 466238 800
rect 470414 0 470470 800
rect 474646 0 474702 800
rect 478878 0 478934 800
rect 483110 0 483166 800
rect 487342 0 487398 800
rect 491574 0 491630 800
rect 495806 0 495862 800
rect 500038 0 500094 800
rect 504270 0 504326 800
rect 508502 0 508558 800
rect 512734 0 512790 800
rect 516966 0 517022 800
rect 521198 0 521254 800
rect 525430 0 525486 800
rect 529662 0 529718 800
rect 533894 0 533950 800
rect 538126 0 538182 800
rect 542358 0 542414 800
rect 546590 0 546646 800
rect 550822 0 550878 800
rect 555054 0 555110 800
<< obsm2 >>
rect 4214 856 557482 349829
rect 4214 546 4838 856
rect 5006 546 9070 856
rect 9238 546 13302 856
rect 13470 546 17534 856
rect 17702 546 21766 856
rect 21934 546 25998 856
rect 26166 546 30230 856
rect 30398 546 34462 856
rect 34630 546 38694 856
rect 38862 546 42926 856
rect 43094 546 47158 856
rect 47326 546 51390 856
rect 51558 546 55622 856
rect 55790 546 59854 856
rect 60022 546 64086 856
rect 64254 546 68318 856
rect 68486 546 72550 856
rect 72718 546 76782 856
rect 76950 546 81014 856
rect 81182 546 85246 856
rect 85414 546 89478 856
rect 89646 546 93710 856
rect 93878 546 97942 856
rect 98110 546 102174 856
rect 102342 546 106406 856
rect 106574 546 110638 856
rect 110806 546 114870 856
rect 115038 546 119102 856
rect 119270 546 123334 856
rect 123502 546 127566 856
rect 127734 546 131798 856
rect 131966 546 136030 856
rect 136198 546 140262 856
rect 140430 546 144494 856
rect 144662 546 148726 856
rect 148894 546 152958 856
rect 153126 546 157190 856
rect 157358 546 161422 856
rect 161590 546 165654 856
rect 165822 546 169886 856
rect 170054 546 174118 856
rect 174286 546 178350 856
rect 178518 546 182582 856
rect 182750 546 186814 856
rect 186982 546 191046 856
rect 191214 546 195278 856
rect 195446 546 199510 856
rect 199678 546 203742 856
rect 203910 546 207974 856
rect 208142 546 212206 856
rect 212374 546 216438 856
rect 216606 546 220670 856
rect 220838 546 224902 856
rect 225070 546 229134 856
rect 229302 546 233366 856
rect 233534 546 237598 856
rect 237766 546 241830 856
rect 241998 546 246062 856
rect 246230 546 250294 856
rect 250462 546 254526 856
rect 254694 546 258758 856
rect 258926 546 262990 856
rect 263158 546 267222 856
rect 267390 546 271454 856
rect 271622 546 275686 856
rect 275854 546 279918 856
rect 280086 546 284150 856
rect 284318 546 288382 856
rect 288550 546 292614 856
rect 292782 546 296846 856
rect 297014 546 301078 856
rect 301246 546 305310 856
rect 305478 546 309542 856
rect 309710 546 313774 856
rect 313942 546 318006 856
rect 318174 546 322238 856
rect 322406 546 326470 856
rect 326638 546 330702 856
rect 330870 546 334934 856
rect 335102 546 339166 856
rect 339334 546 343398 856
rect 343566 546 347630 856
rect 347798 546 351862 856
rect 352030 546 356094 856
rect 356262 546 360326 856
rect 360494 546 364558 856
rect 364726 546 368790 856
rect 368958 546 373022 856
rect 373190 546 377254 856
rect 377422 546 381486 856
rect 381654 546 385718 856
rect 385886 546 389950 856
rect 390118 546 394182 856
rect 394350 546 398414 856
rect 398582 546 402646 856
rect 402814 546 406878 856
rect 407046 546 411110 856
rect 411278 546 415342 856
rect 415510 546 419574 856
rect 419742 546 423806 856
rect 423974 546 428038 856
rect 428206 546 432270 856
rect 432438 546 436502 856
rect 436670 546 440734 856
rect 440902 546 444966 856
rect 445134 546 449198 856
rect 449366 546 453430 856
rect 453598 546 457662 856
rect 457830 546 461894 856
rect 462062 546 466126 856
rect 466294 546 470358 856
rect 470526 546 474590 856
rect 474758 546 478822 856
rect 478990 546 483054 856
rect 483222 546 487286 856
rect 487454 546 491518 856
rect 491686 546 495750 856
rect 495918 546 499982 856
rect 500150 546 504214 856
rect 504382 546 508446 856
rect 508614 546 512678 856
rect 512846 546 516910 856
rect 517078 546 521142 856
rect 521310 546 525374 856
rect 525542 546 529606 856
rect 529774 546 533838 856
rect 534006 546 538070 856
rect 538238 546 542302 856
rect 542470 546 546534 856
rect 546702 546 550766 856
rect 550934 546 554998 856
rect 555166 546 557482 856
<< obsm3 >>
rect 4210 1803 557486 349825
<< metal4 >>
rect 4208 2128 4528 349840
rect 19568 2128 19888 349840
rect 34928 2128 35248 349840
rect 50288 2128 50608 349840
rect 65648 2128 65968 349840
rect 81008 2128 81328 349840
rect 96368 2128 96688 349840
rect 111728 2128 112048 349840
rect 127088 2128 127408 349840
rect 142448 2128 142768 349840
rect 157808 2128 158128 349840
rect 173168 2128 173488 349840
rect 188528 2128 188848 349840
rect 203888 2128 204208 349840
rect 219248 2128 219568 349840
rect 234608 2128 234928 349840
rect 249968 2128 250288 349840
rect 265328 2128 265648 349840
rect 280688 2128 281008 349840
rect 296048 2128 296368 349840
rect 311408 2128 311728 349840
rect 326768 2128 327088 349840
rect 342128 2128 342448 349840
rect 357488 2128 357808 349840
rect 372848 2128 373168 349840
rect 388208 2128 388528 349840
rect 403568 2128 403888 349840
rect 418928 2128 419248 349840
rect 434288 2128 434608 349840
rect 449648 2128 449968 349840
rect 465008 2128 465328 349840
rect 480368 2128 480688 349840
rect 495728 2128 496048 349840
rect 511088 2128 511408 349840
rect 526448 2128 526768 349840
rect 541808 2128 542128 349840
rect 557168 2128 557488 349840
<< labels >>
rlabel metal2 s 26054 0 26110 800 6 ack
port 1 nsew signal output
rlabel metal2 s 186870 0 186926 800 6 adr[0]
port 2 nsew signal input
rlabel metal2 s 229190 0 229246 800 6 adr[10]
port 3 nsew signal input
rlabel metal2 s 233422 0 233478 800 6 adr[11]
port 4 nsew signal input
rlabel metal2 s 237654 0 237710 800 6 adr[12]
port 5 nsew signal input
rlabel metal2 s 241886 0 241942 800 6 adr[13]
port 6 nsew signal input
rlabel metal2 s 246118 0 246174 800 6 adr[14]
port 7 nsew signal input
rlabel metal2 s 250350 0 250406 800 6 adr[15]
port 8 nsew signal input
rlabel metal2 s 254582 0 254638 800 6 adr[16]
port 9 nsew signal input
rlabel metal2 s 258814 0 258870 800 6 adr[17]
port 10 nsew signal input
rlabel metal2 s 263046 0 263102 800 6 adr[18]
port 11 nsew signal input
rlabel metal2 s 267278 0 267334 800 6 adr[19]
port 12 nsew signal input
rlabel metal2 s 191102 0 191158 800 6 adr[1]
port 13 nsew signal input
rlabel metal2 s 271510 0 271566 800 6 adr[20]
port 14 nsew signal input
rlabel metal2 s 275742 0 275798 800 6 adr[21]
port 15 nsew signal input
rlabel metal2 s 279974 0 280030 800 6 adr[22]
port 16 nsew signal input
rlabel metal2 s 284206 0 284262 800 6 adr[23]
port 17 nsew signal input
rlabel metal2 s 288438 0 288494 800 6 adr[24]
port 18 nsew signal input
rlabel metal2 s 292670 0 292726 800 6 adr[25]
port 19 nsew signal input
rlabel metal2 s 296902 0 296958 800 6 adr[26]
port 20 nsew signal input
rlabel metal2 s 301134 0 301190 800 6 adr[27]
port 21 nsew signal input
rlabel metal2 s 305366 0 305422 800 6 adr[28]
port 22 nsew signal input
rlabel metal2 s 309598 0 309654 800 6 adr[29]
port 23 nsew signal input
rlabel metal2 s 195334 0 195390 800 6 adr[2]
port 24 nsew signal input
rlabel metal2 s 313830 0 313886 800 6 adr[30]
port 25 nsew signal input
rlabel metal2 s 318062 0 318118 800 6 adr[31]
port 26 nsew signal input
rlabel metal2 s 199566 0 199622 800 6 adr[3]
port 27 nsew signal input
rlabel metal2 s 203798 0 203854 800 6 adr[4]
port 28 nsew signal input
rlabel metal2 s 208030 0 208086 800 6 adr[5]
port 29 nsew signal input
rlabel metal2 s 212262 0 212318 800 6 adr[6]
port 30 nsew signal input
rlabel metal2 s 216494 0 216550 800 6 adr[7]
port 31 nsew signal input
rlabel metal2 s 220726 0 220782 800 6 adr[8]
port 32 nsew signal input
rlabel metal2 s 224958 0 225014 800 6 adr[9]
port 33 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 clk
port 34 nsew signal input
rlabel metal2 s 508502 0 508558 800 6 column[0]
port 35 nsew signal output
rlabel metal2 s 550822 0 550878 800 6 column[10]
port 36 nsew signal output
rlabel metal2 s 555054 0 555110 800 6 column[11]
port 37 nsew signal output
rlabel metal2 s 512734 0 512790 800 6 column[1]
port 38 nsew signal output
rlabel metal2 s 516966 0 517022 800 6 column[2]
port 39 nsew signal output
rlabel metal2 s 521198 0 521254 800 6 column[3]
port 40 nsew signal output
rlabel metal2 s 525430 0 525486 800 6 column[4]
port 41 nsew signal output
rlabel metal2 s 529662 0 529718 800 6 column[5]
port 42 nsew signal output
rlabel metal2 s 533894 0 533950 800 6 column[6]
port 43 nsew signal output
rlabel metal2 s 538126 0 538182 800 6 column[7]
port 44 nsew signal output
rlabel metal2 s 542358 0 542414 800 6 column[8]
port 45 nsew signal output
rlabel metal2 s 546590 0 546646 800 6 column[9]
port 46 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 cyc
port 47 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 dat[0]
port 48 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 dat[10]
port 49 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 dat[11]
port 50 nsew signal input
rlabel metal2 s 102230 0 102286 800 6 dat[12]
port 51 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 dat[13]
port 52 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 dat[14]
port 53 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 dat[15]
port 54 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 dat[16]
port 55 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 dat[17]
port 56 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 dat[18]
port 57 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 dat[19]
port 58 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 dat[1]
port 59 nsew signal input
rlabel metal2 s 136086 0 136142 800 6 dat[20]
port 60 nsew signal input
rlabel metal2 s 140318 0 140374 800 6 dat[21]
port 61 nsew signal input
rlabel metal2 s 144550 0 144606 800 6 dat[22]
port 62 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 dat[23]
port 63 nsew signal input
rlabel metal2 s 153014 0 153070 800 6 dat[24]
port 64 nsew signal input
rlabel metal2 s 157246 0 157302 800 6 dat[25]
port 65 nsew signal input
rlabel metal2 s 161478 0 161534 800 6 dat[26]
port 66 nsew signal input
rlabel metal2 s 165710 0 165766 800 6 dat[27]
port 67 nsew signal input
rlabel metal2 s 169942 0 169998 800 6 dat[28]
port 68 nsew signal input
rlabel metal2 s 174174 0 174230 800 6 dat[29]
port 69 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 dat[2]
port 70 nsew signal input
rlabel metal2 s 178406 0 178462 800 6 dat[30]
port 71 nsew signal input
rlabel metal2 s 182638 0 182694 800 6 dat[31]
port 72 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 dat[3]
port 73 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 dat[4]
port 74 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 dat[5]
port 75 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 dat[6]
port 76 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 dat[7]
port 77 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 dat[8]
port 78 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 dat[9]
port 79 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 display_enable
port 80 nsew signal output
rlabel metal2 s 322294 0 322350 800 6 dout[0]
port 81 nsew signal output
rlabel metal2 s 364614 0 364670 800 6 dout[10]
port 82 nsew signal output
rlabel metal2 s 368846 0 368902 800 6 dout[11]
port 83 nsew signal output
rlabel metal2 s 373078 0 373134 800 6 dout[12]
port 84 nsew signal output
rlabel metal2 s 377310 0 377366 800 6 dout[13]
port 85 nsew signal output
rlabel metal2 s 381542 0 381598 800 6 dout[14]
port 86 nsew signal output
rlabel metal2 s 385774 0 385830 800 6 dout[15]
port 87 nsew signal output
rlabel metal2 s 390006 0 390062 800 6 dout[16]
port 88 nsew signal output
rlabel metal2 s 394238 0 394294 800 6 dout[17]
port 89 nsew signal output
rlabel metal2 s 398470 0 398526 800 6 dout[18]
port 90 nsew signal output
rlabel metal2 s 402702 0 402758 800 6 dout[19]
port 91 nsew signal output
rlabel metal2 s 326526 0 326582 800 6 dout[1]
port 92 nsew signal output
rlabel metal2 s 406934 0 406990 800 6 dout[20]
port 93 nsew signal output
rlabel metal2 s 411166 0 411222 800 6 dout[21]
port 94 nsew signal output
rlabel metal2 s 415398 0 415454 800 6 dout[22]
port 95 nsew signal output
rlabel metal2 s 419630 0 419686 800 6 dout[23]
port 96 nsew signal output
rlabel metal2 s 423862 0 423918 800 6 dout[24]
port 97 nsew signal output
rlabel metal2 s 428094 0 428150 800 6 dout[25]
port 98 nsew signal output
rlabel metal2 s 432326 0 432382 800 6 dout[26]
port 99 nsew signal output
rlabel metal2 s 436558 0 436614 800 6 dout[27]
port 100 nsew signal output
rlabel metal2 s 440790 0 440846 800 6 dout[28]
port 101 nsew signal output
rlabel metal2 s 445022 0 445078 800 6 dout[29]
port 102 nsew signal output
rlabel metal2 s 330758 0 330814 800 6 dout[2]
port 103 nsew signal output
rlabel metal2 s 449254 0 449310 800 6 dout[30]
port 104 nsew signal output
rlabel metal2 s 453486 0 453542 800 6 dout[31]
port 105 nsew signal output
rlabel metal2 s 334990 0 335046 800 6 dout[3]
port 106 nsew signal output
rlabel metal2 s 339222 0 339278 800 6 dout[4]
port 107 nsew signal output
rlabel metal2 s 343454 0 343510 800 6 dout[5]
port 108 nsew signal output
rlabel metal2 s 347686 0 347742 800 6 dout[6]
port 109 nsew signal output
rlabel metal2 s 351918 0 351974 800 6 dout[7]
port 110 nsew signal output
rlabel metal2 s 356150 0 356206 800 6 dout[8]
port 111 nsew signal output
rlabel metal2 s 360382 0 360438 800 6 dout[9]
port 112 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 h_sync
port 113 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 n_blank
port 114 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 n_sync
port 115 nsew signal output
rlabel metal2 s 457718 0 457774 800 6 row[0]
port 116 nsew signal output
rlabel metal2 s 500038 0 500094 800 6 row[10]
port 117 nsew signal output
rlabel metal2 s 504270 0 504326 800 6 row[11]
port 118 nsew signal output
rlabel metal2 s 461950 0 462006 800 6 row[1]
port 119 nsew signal output
rlabel metal2 s 466182 0 466238 800 6 row[2]
port 120 nsew signal output
rlabel metal2 s 470414 0 470470 800 6 row[3]
port 121 nsew signal output
rlabel metal2 s 474646 0 474702 800 6 row[4]
port 122 nsew signal output
rlabel metal2 s 478878 0 478934 800 6 row[5]
port 123 nsew signal output
rlabel metal2 s 483110 0 483166 800 6 row[6]
port 124 nsew signal output
rlabel metal2 s 487342 0 487398 800 6 row[7]
port 125 nsew signal output
rlabel metal2 s 491574 0 491630 800 6 row[8]
port 126 nsew signal output
rlabel metal2 s 495806 0 495862 800 6 row[9]
port 127 nsew signal output
rlabel metal2 s 9126 0 9182 800 6 rst
port 128 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 stb
port 129 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 v_sync
port 130 nsew signal output
rlabel metal4 s 4208 2128 4528 349840 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 349840 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 349840 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 349840 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 349840 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 349840 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 349840 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 349840 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 349840 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 349840 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 349840 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 349840 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 349840 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 349840 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 349840 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 349840 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 349840 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 349840 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 557168 2128 557488 349840 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 349840 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 349840 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 349840 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 349840 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 349840 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 349840 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 349840 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 349840 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 349840 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 349840 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 349840 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 349840 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 349840 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 349840 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 349840 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 349840 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 349840 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 541808 2128 542128 349840 6 vssd1
port 132 nsew ground bidirectional
rlabel metal2 s 21822 0 21878 800 6 we
port 133 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 560000 352000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 52885636
string GDS_FILE /home/m/Wishbone_VGA_controller/openlane/Wishbone_VGA_controller/runs/23_06_03_18_22/results/signoff/Wishbone_VGA_controller.magic.gds
string GDS_START 808916
<< end >>

