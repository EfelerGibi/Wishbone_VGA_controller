magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< locali >>
rect 11923 32808 11954 32846
rect 18056 32815 18086 32844
rect 18234 32813 18269 32838
rect 18234 32803 18242 32813
rect 16799 32751 16831 32795
rect 16965 32758 16996 32798
rect 18216 32779 18242 32781
rect 18420 32797 18456 32833
rect 18276 32779 18282 32781
rect 18216 32741 18282 32779
rect 19211 32744 19267 32788
rect 18216 32707 18242 32741
rect 18276 32707 18282 32741
<< viali >>
rect 18242 32779 18276 32813
rect 18242 32707 18276 32741
<< metal1 >>
rect 18522 33471 19108 33673
rect 17266 33331 17272 33383
rect 17324 33331 17336 33383
rect 17388 33331 17394 33383
rect 17875 33269 18003 33399
tri 27460 33067 27488 33095 ne
rect 18228 32814 18282 32825
rect 18280 32762 18282 32814
rect 18228 32750 18282 32762
rect 18280 32698 18282 32750
rect 18228 32692 18282 32698
rect 11513 32365 11551 32404
rect 18581 32317 19176 32472
tri 27665 32197 27695 32227 ne
rect 27695 32197 27698 32227
rect 27140 32164 27192 32197
tri 27695 32194 27698 32197 ne
tri 27750 32194 27783 32227 nw
rect 19853 31506 19905 31512
rect 19853 31442 19905 31454
rect 19853 31384 19905 31390
rect 24432 30637 24634 30679
rect 25923 30641 26053 30683
rect 26335 30641 26537 30683
rect 26861 30641 27063 30683
rect 27575 30646 27721 30683
rect 27321 30418 27352 30562
tri 26781 29926 26787 29932 se
rect 26787 29926 26833 30165
rect 26781 29920 26833 29926
tri 27359 29893 27365 29899 nw
rect 26781 29856 26833 29868
rect 26781 29798 26833 29804
rect 24184 29706 24386 29748
rect 27091 24877 27137 24917
rect 27091 24740 27137 24781
rect 26721 23039 26752 23133
rect 27171 22975 27217 23015
rect 27289 22777 27335 22823
rect 26650 22321 26674 22407
rect 27289 21535 27335 21581
rect 25465 20856 25511 20902
rect 27247 20545 27293 20585
rect 25923 17881 26053 17923
rect 26335 17905 26537 17947
rect 24184 17775 24386 17817
rect 24710 17775 24912 17817
rect 25307 17775 25437 17817
rect 26861 17775 27063 17817
rect 27575 17775 27721 17812
<< via1 >>
rect 17272 33331 17324 33383
rect 17336 33331 17388 33383
rect 18228 32813 18280 32814
rect 18228 32779 18242 32813
rect 18242 32779 18276 32813
rect 18276 32779 18280 32813
rect 18228 32762 18280 32779
rect 18228 32741 18280 32750
rect 18228 32707 18242 32741
rect 18242 32707 18276 32741
rect 18276 32707 18280 32741
rect 18228 32698 18280 32707
rect 19853 31454 19905 31506
rect 19853 31390 19905 31442
rect 26781 29868 26833 29920
rect 26781 29804 26833 29856
<< metal2 >>
rect 11274 33500 11643 33685
rect 17260 33453 17269 33509
rect 17325 33453 17349 33509
rect 17405 33453 17414 33509
rect 17266 33383 17394 33453
tri 17394 33433 17414 33453 nw
rect 17266 33331 17272 33383
rect 17324 33331 17336 33383
rect 17388 33331 17394 33383
rect 20036 33327 20045 33383
rect 20101 33327 20125 33383
rect 20181 33327 20190 33383
tri 20037 33322 20042 33327 ne
rect 20042 33322 20127 33327
tri 20127 33322 20132 33327 nw
tri 15704 33201 15760 33257 se
rect 15760 33201 16206 33257
rect 16262 33201 16307 33257
rect 16363 33201 16408 33257
rect 16464 33201 16473 33257
tri 15658 33155 15704 33201 se
rect 15704 33155 15736 33201
tri 15736 33155 15782 33201 nw
tri 15580 33077 15658 33155 se
tri 15658 33077 15736 33155 nw
tri 15811 33077 15865 33131 se
rect 15865 33077 16206 33131
tri 15502 32999 15580 33077 se
tri 15580 32999 15658 33077 nw
tri 15787 33053 15811 33077 se
rect 15811 33075 16206 33077
rect 16262 33075 16307 33131
rect 16363 33075 16408 33131
rect 16464 33075 16473 33131
rect 15811 33053 15865 33075
tri 15865 33053 15887 33075 nw
tri 15733 32999 15787 33053 se
tri 15424 32921 15502 32999 se
tri 15502 32921 15580 32999 nw
tri 15709 32975 15733 32999 se
rect 15733 32975 15787 32999
tri 15787 32975 15865 33053 nw
tri 15655 32921 15709 32975 se
tri 15402 32899 15424 32921 se
rect 14766 32843 14775 32899
rect 14831 32843 14876 32899
rect 14932 32843 14977 32899
rect 15033 32843 15424 32899
tri 15424 32843 15502 32921 nw
tri 15631 32897 15655 32921 se
rect 15655 32897 15709 32921
tri 15709 32897 15787 32975 nw
tri 15577 32843 15631 32897 se
tri 15553 32819 15577 32843 se
rect 15577 32819 15631 32843
tri 15631 32819 15709 32897 nw
rect 16933 32823 16942 32879
rect 16998 32823 17022 32879
rect 17078 32823 17087 32879
tri 15548 32814 15553 32819 se
rect 15553 32814 15626 32819
tri 15626 32814 15631 32819 nw
tri 15507 32773 15548 32814 se
rect 15548 32773 15585 32814
tri 15585 32773 15626 32814 nw
rect 16951 32805 17003 32823
rect 18228 32814 18280 32820
rect 14766 32717 14775 32773
rect 14831 32717 14876 32773
rect 14932 32717 14977 32773
rect 15033 32762 15574 32773
tri 15574 32762 15585 32773 nw
rect 15033 32750 15562 32762
tri 15562 32750 15574 32762 nw
rect 18228 32753 18280 32762
rect 15033 32717 15529 32750
tri 15529 32717 15562 32750 nw
rect 18129 32697 18138 32753
rect 18194 32697 18218 32753
rect 18274 32750 18283 32753
rect 18280 32698 18283 32750
rect 18274 32697 18283 32698
rect 18228 32692 18280 32697
tri 19968 31516 20042 31590 se
rect 20042 31516 20097 33322
tri 20097 33292 20127 33322 nw
rect 19853 31506 20097 31516
rect 19905 31454 20097 31506
rect 19853 31442 20097 31454
rect 19905 31390 20097 31442
rect 19853 31384 20097 31390
rect 24402 29926 24458 29929
tri 24458 29926 24461 29929 sw
rect 24402 29920 26833 29926
tri 23413 29868 23418 29873 sw
rect 23413 29856 23418 29868
tri 23418 29856 23430 29868 sw
rect 24458 29868 26781 29920
rect 24458 29864 26833 29868
rect 24402 29856 26833 29864
rect 23413 29842 23430 29856
tri 23430 29842 23444 29856 sw
rect 24402 29840 26781 29856
tri 23409 29775 23419 29785 ne
rect 23419 29775 23443 29785
rect 24458 29804 26781 29840
rect 24458 29798 26833 29804
rect 24402 29775 24458 29784
tri 24458 29775 24481 29798 nw
tri 23419 29751 23443 29775 ne
rect 2214 29431 2333 29489
rect 5497 29432 5506 29488
rect 5562 29432 5586 29488
rect 5642 29432 5651 29488
rect 2028 29282 2200 29364
rect 5291 29332 5300 29388
rect 5356 29332 5380 29388
rect 5436 29332 5445 29388
rect 4839 28595 4994 28884
rect 18919 27043 19027 27411
rect 22701 27039 22809 27407
rect 26693 23756 26745 23808
rect 25722 23272 25873 23315
rect 25032 21231 25088 21240
rect 25032 21151 25088 21175
rect 25032 21086 25088 21095
rect 25159 21137 25465 21146
rect 25215 21081 25465 21137
rect 25159 21057 25465 21081
rect 25215 21018 25465 21057
rect 25159 20992 25215 21001
rect 24780 20822 24836 20831
rect 25098 20781 25150 20828
rect 24780 20742 24836 20766
rect 24780 20677 24836 20686
rect 26781 20301 26833 20359
tri 27553 20199 27585 20231 ne
rect 24906 20105 24962 20114
tri 24962 20081 24995 20114 sw
rect 24962 20076 26751 20081
tri 26751 20076 26756 20081 sw
rect 24962 20064 26756 20076
tri 26756 20064 26768 20076 sw
tri 27573 20064 27585 20076 se
rect 27585 20064 27671 20231
tri 27671 20199 27703 20231 nw
rect 24962 20049 26768 20064
rect 24906 20025 26768 20049
rect 24962 19995 26768 20025
tri 26768 19995 26837 20064 sw
tri 27504 19995 27573 20064 se
rect 27573 20040 27671 20064
rect 27573 19995 27585 20040
rect 24906 19960 24962 19969
tri 24962 19961 24996 19995 nw
tri 26715 19961 26749 19995 ne
rect 26749 19961 26837 19995
tri 26837 19961 26871 19995 sw
tri 27470 19961 27504 19995 se
rect 27504 19961 27585 19995
tri 26749 19960 26750 19961 ne
rect 26750 19960 26871 19961
tri 26750 19942 26768 19960 ne
rect 26768 19954 26871 19960
tri 26871 19954 26878 19961 sw
tri 27463 19954 27470 19961 se
rect 27470 19954 27585 19961
tri 27585 19954 27671 20040 nw
rect 26768 19942 26878 19954
tri 26878 19942 26890 19954 sw
tri 27451 19942 27463 19954 se
rect 27463 19942 27573 19954
tri 27573 19942 27585 19954 nw
tri 26768 19856 26854 19942 ne
rect 26854 19856 27487 19942
tri 27487 19856 27573 19942 nw
tri 24648 18592 24654 18598 se
rect 24654 18592 24710 18598
tri 24710 18592 24716 18598 sw
tri 24644 18588 24648 18592 se
rect 24648 18589 24716 18592
rect 24648 18588 24654 18589
rect 24710 18588 24716 18589
tri 24716 18588 24720 18592 sw
tri 25406 18588 25410 18592 se
rect 25410 18588 25468 18592
tri 25468 18588 25472 18592 sw
rect 24654 18509 24710 18533
tri 24638 18444 24654 18460 ne
tri 25376 18460 25388 18472 ne
rect 25388 18460 25410 18472
rect 24654 18444 24710 18453
tri 24710 18444 24726 18460 nw
tri 25388 18444 25404 18460 ne
rect 25404 18444 25410 18460
tri 25404 18438 25410 18444 ne
tri 25466 18438 25500 18472 nw
rect 26621 17940 26673 17987
<< via2 >>
rect 17269 33453 17325 33509
rect 17349 33453 17405 33509
rect 20045 33327 20101 33383
rect 20125 33327 20181 33383
rect 16206 33201 16262 33257
rect 16307 33201 16363 33257
rect 16408 33201 16464 33257
rect 16206 33075 16262 33131
rect 16307 33075 16363 33131
rect 16408 33075 16464 33131
rect 14775 32843 14831 32899
rect 14876 32843 14932 32899
rect 14977 32843 15033 32899
rect 16942 32823 16998 32879
rect 17022 32823 17078 32879
rect 14775 32717 14831 32773
rect 14876 32717 14932 32773
rect 14977 32717 15033 32773
rect 18138 32697 18194 32753
rect 18218 32750 18274 32753
rect 18218 32698 18228 32750
rect 18228 32698 18274 32750
rect 18218 32697 18274 32698
rect 24402 29864 24458 29920
rect 24402 29784 24458 29840
rect 5506 29432 5562 29488
rect 5586 29432 5642 29488
rect 5300 29332 5356 29388
rect 5380 29332 5436 29388
rect 25032 21175 25088 21231
rect 25032 21095 25088 21151
rect 25159 21081 25215 21137
rect 25159 21001 25215 21057
rect 24780 20766 24836 20822
rect 24780 20686 24836 20742
rect 24906 20049 24962 20105
rect 24906 19969 24962 20025
rect 24654 18533 24710 18589
rect 24654 18453 24710 18509
<< metal3 >>
rect 17264 33509 23690 33514
rect 17264 33453 17269 33509
rect 17325 33453 17349 33509
rect 17405 33488 23690 33509
tri 23690 33488 23716 33514 sw
rect 17405 33453 23716 33488
rect 17264 33448 23716 33453
tri 23662 33394 23716 33448 ne
tri 23716 33394 23810 33488 sw
tri 23716 33388 23722 33394 ne
rect 23722 33388 23810 33394
tri 23810 33388 23816 33394 sw
rect 20040 33383 23635 33388
rect 20040 33327 20045 33383
rect 20101 33327 20125 33383
rect 20181 33340 23635 33383
tri 23635 33340 23683 33388 sw
tri 23722 33340 23770 33388 ne
rect 23770 33340 23816 33388
tri 23816 33340 23864 33388 sw
rect 20181 33327 23683 33340
rect 20040 33322 23683 33327
tri 23683 33322 23701 33340 sw
tri 23770 33322 23788 33340 ne
rect 23788 33322 23864 33340
tri 23864 33322 23882 33340 sw
tri 23607 33262 23667 33322 ne
rect 23667 33307 23701 33322
tri 23701 33307 23716 33322 sw
tri 23788 33307 23803 33322 ne
rect 23803 33307 23882 33322
rect 23667 33300 23716 33307
tri 23716 33300 23723 33307 sw
tri 23803 33300 23810 33307 ne
rect 23810 33300 23882 33307
tri 23882 33300 23904 33322 sw
rect 23667 33262 23723 33300
tri 23723 33262 23761 33300 sw
tri 23810 33262 23848 33300 ne
rect 23848 33262 23904 33300
tri 23904 33262 23942 33300 sw
rect 16183 33257 23581 33262
rect 16183 33201 16206 33257
rect 16262 33201 16307 33257
rect 16363 33201 16408 33257
rect 16464 33246 23581 33257
tri 23581 33246 23597 33262 sw
tri 23667 33246 23683 33262 ne
rect 23683 33246 23761 33262
tri 23761 33246 23777 33262 sw
tri 23848 33246 23864 33262 ne
rect 23864 33246 23942 33262
tri 23942 33246 23958 33262 sw
rect 16464 33201 23597 33246
rect 16183 33196 23597 33201
tri 23597 33196 23647 33246 sw
tri 23683 33196 23733 33246 ne
rect 23733 33213 23777 33246
tri 23777 33213 23810 33246 sw
tri 23864 33213 23897 33246 ne
rect 23897 33213 23958 33246
rect 23733 33206 23810 33213
tri 23810 33206 23817 33213 sw
tri 23897 33206 23904 33213 ne
rect 23904 33206 23958 33213
tri 23958 33206 23998 33246 sw
rect 23733 33196 23817 33206
tri 23817 33196 23827 33206 sw
tri 23904 33196 23914 33206 ne
rect 23914 33196 23998 33206
tri 23998 33196 24008 33206 sw
tri 23553 33192 23557 33196 ne
rect 23557 33192 23647 33196
tri 23647 33192 23651 33196 sw
tri 23733 33192 23737 33196 ne
rect 23737 33192 23827 33196
tri 23557 33168 23581 33192 ne
rect 23581 33184 23651 33192
tri 23651 33184 23659 33192 sw
tri 23737 33184 23745 33192 ne
rect 23745 33184 23827 33192
rect 23581 33168 23659 33184
tri 23581 33136 23613 33168 ne
rect 23613 33152 23659 33168
tri 23659 33152 23691 33184 sw
tri 23745 33152 23777 33184 ne
rect 23777 33152 23827 33184
tri 23827 33152 23871 33196 sw
tri 23914 33152 23958 33196 ne
rect 23958 33152 24008 33196
tri 24008 33152 24052 33196 sw
rect 23613 33136 23691 33152
tri 23691 33136 23707 33152 sw
tri 23777 33136 23793 33152 ne
rect 23793 33136 23871 33152
tri 23871 33136 23887 33152 sw
tri 23958 33136 23974 33152 ne
rect 23974 33136 24052 33152
tri 24052 33136 24068 33152 sw
rect 16183 33131 23527 33136
rect 16183 33075 16206 33131
rect 16262 33075 16307 33131
rect 16363 33075 16408 33131
rect 16464 33130 23527 33131
tri 23527 33130 23533 33136 sw
tri 23613 33130 23619 33136 ne
rect 23619 33130 23707 33136
rect 16464 33098 23533 33130
tri 23533 33098 23565 33130 sw
tri 23619 33098 23651 33130 ne
rect 23651 33098 23707 33130
tri 23707 33098 23745 33136 sw
tri 23793 33098 23831 33136 ne
rect 23831 33119 23887 33136
tri 23887 33119 23904 33136 sw
tri 23974 33119 23991 33136 ne
rect 23991 33119 24068 33136
rect 23831 33112 23904 33119
tri 23904 33112 23911 33119 sw
tri 23991 33112 23998 33119 ne
rect 23998 33112 24068 33119
tri 24068 33112 24092 33136 sw
rect 23831 33098 23911 33112
rect 16464 33075 23565 33098
rect 16183 33070 23565 33075
tri 23565 33070 23593 33098 sw
tri 23651 33070 23679 33098 ne
rect 23679 33090 23745 33098
tri 23745 33090 23753 33098 sw
tri 23831 33090 23839 33098 ne
rect 23839 33090 23911 33098
rect 23679 33070 23753 33090
tri 23753 33070 23773 33090 sw
tri 23839 33070 23859 33090 ne
rect 23859 33070 23911 33090
tri 23911 33070 23953 33112 sw
tri 23998 33070 24040 33112 ne
rect 24040 33070 24092 33112
tri 24092 33070 24134 33112 sw
tri 23499 33044 23525 33070 ne
rect 23525 33044 23593 33070
tri 23593 33044 23619 33070 sw
tri 23679 33044 23705 33070 ne
rect 23705 33058 23773 33070
tri 23773 33058 23785 33070 sw
tri 23859 33058 23871 33070 ne
rect 23871 33058 23953 33070
tri 23953 33058 23965 33070 sw
tri 24040 33058 24052 33070 ne
rect 24052 33058 24134 33070
tri 24134 33058 24146 33070 sw
rect 23705 33044 23785 33058
tri 23525 33042 23527 33044 ne
rect 23527 33042 23619 33044
tri 23527 33010 23559 33042 ne
rect 23559 33036 23619 33042
tri 23619 33036 23627 33044 sw
tri 23705 33036 23713 33044 ne
rect 23713 33036 23785 33044
rect 23559 33010 23627 33036
tri 23627 33010 23653 33036 sw
tri 23713 33010 23739 33036 ne
rect 23739 33010 23785 33036
tri 23785 33010 23833 33058 sw
tri 23871 33010 23919 33058 ne
rect 23919 33025 23965 33058
tri 23965 33025 23998 33058 sw
tri 24052 33025 24085 33058 ne
rect 24085 33025 24146 33058
rect 23919 33018 23998 33025
tri 23998 33018 24005 33025 sw
tri 24085 33018 24092 33025 ne
rect 24092 33018 24146 33025
tri 24146 33018 24186 33058 sw
rect 23919 33010 24005 33018
tri 24005 33010 24013 33018 sw
tri 24092 33010 24100 33018 ne
rect 24100 33010 24186 33018
tri 24186 33010 24194 33018 sw
rect 16649 32990 23473 33010
tri 23473 32990 23493 33010 sw
tri 23559 32990 23579 33010 ne
rect 23579 33004 23653 33010
tri 23653 33004 23659 33010 sw
tri 23739 33004 23745 33010 ne
rect 23745 33004 23833 33010
tri 23833 33004 23839 33010 sw
tri 23919 33004 23925 33010 ne
rect 23925 33004 24013 33010
rect 23579 32990 23659 33004
tri 23659 32990 23673 33004 sw
tri 23745 32990 23759 33004 ne
rect 23759 32996 23839 33004
tri 23839 32996 23847 33004 sw
tri 23925 32996 23933 33004 ne
rect 23933 32996 24013 33004
rect 23759 32990 23847 32996
tri 23847 32990 23853 32996 sw
tri 23933 32990 23939 32996 ne
rect 23939 32990 24013 32996
tri 24013 32990 24033 33010 sw
tri 24100 32990 24120 33010 ne
rect 24120 32990 24194 33010
tri 24194 32990 24214 33010 sw
rect 16649 32956 23493 32990
tri 23493 32956 23527 32990 sw
tri 23579 32956 23613 32990 ne
rect 23613 32956 23673 32990
rect 16649 32950 23527 32956
tri 23527 32950 23533 32956 sw
tri 23613 32950 23619 32956 ne
rect 23619 32950 23673 32956
tri 23673 32950 23713 32990 sw
tri 23759 32950 23799 32990 ne
rect 23799 32964 23853 32990
tri 23853 32964 23879 32990 sw
tri 23939 32964 23965 32990 ne
rect 23965 32964 24033 32990
tri 24033 32964 24059 32990 sw
tri 24120 32964 24146 32990 ne
rect 24146 32964 24214 32990
tri 24214 32964 24240 32990 sw
rect 23799 32950 23879 32964
rect 16649 32944 23533 32950
tri 23445 32904 23485 32944 ne
rect 23485 32904 23533 32944
tri 23533 32904 23579 32950 sw
tri 23619 32904 23665 32950 ne
rect 23665 32942 23713 32950
tri 23713 32942 23721 32950 sw
tri 23799 32942 23807 32950 ne
rect 23807 32942 23879 32950
rect 23665 32910 23721 32942
tri 23721 32910 23753 32942 sw
tri 23807 32910 23839 32942 ne
rect 23839 32910 23879 32942
tri 23879 32910 23933 32964 sw
tri 23965 32910 24019 32964 ne
rect 24019 32931 24059 32964
tri 24059 32931 24092 32964 sw
tri 24146 32931 24179 32964 ne
rect 24179 32931 24240 32964
rect 24019 32924 24092 32931
tri 24092 32924 24099 32931 sw
tri 24179 32924 24186 32931 ne
rect 24186 32924 24240 32931
tri 24240 32924 24280 32964 sw
rect 24019 32910 24099 32924
rect 23665 32904 23753 32910
tri 23753 32904 23759 32910 sw
tri 23839 32904 23845 32910 ne
rect 23845 32904 23933 32910
tri 23933 32904 23939 32910 sw
tri 24019 32904 24025 32910 ne
rect 24025 32904 24099 32910
tri 24099 32904 24119 32924 sw
tri 24186 32904 24206 32924 ne
rect 24206 32904 24280 32924
tri 24280 32904 24300 32924 sw
tri 5608 32899 5613 32904 se
rect 5613 32899 15041 32904
tri 5593 32884 5608 32899 se
rect 5608 32884 14775 32899
tri 5552 32843 5593 32884 se
rect 5593 32843 14775 32884
rect 14831 32843 14876 32899
rect 14932 32843 14977 32899
rect 15033 32843 15041 32899
tri 23485 32896 23493 32904 ne
rect 23493 32896 23579 32904
tri 23579 32896 23587 32904 sw
tri 23665 32896 23673 32904 ne
rect 23673 32896 23759 32904
tri 23759 32896 23767 32904 sw
tri 23845 32896 23853 32904 ne
rect 23853 32902 23939 32904
tri 23939 32902 23941 32904 sw
tri 24025 32902 24027 32904 ne
rect 24027 32902 24119 32904
rect 23853 32896 23941 32902
tri 23941 32896 23947 32902 sw
tri 24027 32896 24033 32902 ne
rect 24033 32896 24119 32902
tri 24119 32896 24127 32904 sw
tri 24206 32896 24214 32904 ne
rect 24214 32896 24300 32904
tri 24300 32896 24308 32904 sw
tri 23493 32884 23505 32896 ne
rect 23505 32884 23587 32896
tri 23587 32884 23599 32896 sw
tri 23673 32884 23685 32896 ne
rect 23685 32884 23767 32896
tri 23767 32884 23779 32896 sw
tri 23853 32884 23865 32896 ne
rect 23865 32884 23947 32896
tri 23947 32884 23959 32896 sw
tri 24033 32884 24045 32896 ne
rect 24045 32884 24127 32896
tri 24127 32884 24139 32896 sw
tri 24214 32884 24226 32896 ne
rect 24226 32884 24308 32896
tri 24308 32884 24320 32896 sw
tri 5532 32823 5552 32843 se
rect 5552 32838 15041 32843
rect 16937 32879 23419 32884
rect 5552 32823 5660 32838
tri 5660 32823 5675 32838 nw
rect 16937 32823 16942 32879
rect 16998 32823 17022 32879
rect 17078 32842 23419 32879
tri 23419 32842 23461 32884 sw
tri 23505 32842 23547 32884 ne
rect 23547 32864 23599 32884
tri 23599 32864 23619 32884 sw
tri 23685 32864 23705 32884 ne
rect 23705 32864 23779 32884
rect 23547 32856 23619 32864
tri 23619 32856 23627 32864 sw
tri 23705 32856 23713 32864 ne
rect 23713 32856 23779 32864
tri 23779 32856 23807 32884 sw
tri 23865 32856 23893 32884 ne
rect 23893 32870 23959 32884
tri 23959 32870 23973 32884 sw
tri 24045 32870 24059 32884 ne
rect 24059 32870 24139 32884
tri 24139 32870 24153 32884 sw
tri 24226 32870 24240 32884 ne
rect 24240 32870 24320 32884
tri 24320 32870 24334 32884 sw
rect 23893 32856 23973 32870
rect 23547 32842 23627 32856
tri 23627 32842 23641 32856 sw
tri 23713 32842 23727 32856 ne
rect 23727 32848 23807 32856
tri 23807 32848 23815 32856 sw
tri 23893 32848 23901 32856 ne
rect 23901 32848 23973 32856
rect 23727 32842 23815 32848
tri 23815 32842 23821 32848 sw
tri 23901 32842 23907 32848 ne
rect 23907 32842 23973 32848
tri 23973 32842 24001 32870 sw
tri 24059 32842 24087 32870 ne
rect 24087 32842 24153 32870
tri 24153 32842 24181 32870 sw
tri 24240 32842 24268 32870 ne
rect 24268 32842 24334 32870
tri 24334 32842 24362 32870 sw
rect 17078 32823 23461 32842
tri 5527 32818 5532 32823 se
rect 5532 32818 5655 32823
tri 5655 32818 5660 32823 nw
rect 16937 32818 23461 32823
tri 5485 32776 5527 32818 se
rect 5527 32778 5615 32818
tri 5615 32778 5655 32818 nw
tri 23391 32778 23431 32818 ne
rect 23431 32810 23461 32818
tri 23461 32810 23493 32842 sw
tri 23547 32810 23579 32842 ne
rect 23579 32810 23641 32842
rect 23431 32802 23493 32810
tri 23493 32802 23501 32810 sw
tri 23579 32802 23587 32810 ne
rect 23587 32802 23641 32810
tri 23641 32802 23681 32842 sw
tri 23727 32802 23767 32842 ne
rect 23767 32816 23821 32842
tri 23821 32816 23847 32842 sw
tri 23907 32816 23933 32842 ne
rect 23933 32816 24001 32842
tri 24001 32816 24027 32842 sw
tri 24087 32816 24113 32842 ne
rect 24113 32837 24181 32842
tri 24181 32837 24186 32842 sw
tri 24268 32837 24273 32842 ne
rect 24273 32837 24362 32842
rect 24113 32830 24186 32837
tri 24186 32830 24193 32837 sw
tri 24273 32830 24280 32837 ne
rect 24280 32830 24362 32837
tri 24362 32830 24374 32842 sw
rect 24113 32816 24193 32830
rect 23767 32802 23847 32816
tri 23847 32802 23861 32816 sw
tri 23933 32802 23947 32816 ne
rect 23947 32808 24027 32816
tri 24027 32808 24035 32816 sw
tri 24113 32808 24121 32816 ne
rect 24121 32808 24193 32816
rect 23947 32802 24035 32808
tri 24035 32802 24041 32808 sw
tri 24121 32802 24127 32808 ne
rect 24127 32802 24193 32808
tri 24193 32802 24221 32830 sw
tri 24280 32802 24308 32830 ne
rect 24308 32802 24374 32830
tri 24374 32802 24402 32830 sw
rect 23431 32778 23501 32802
rect 5527 32776 5613 32778
tri 5613 32776 5615 32778 nw
tri 5747 32776 5749 32778 se
rect 5749 32776 15041 32778
tri 5482 32773 5485 32776 se
rect 5485 32773 5610 32776
tri 5610 32773 5613 32776 nw
tri 5744 32773 5747 32776 se
rect 5747 32773 15041 32776
tri 5467 32758 5482 32773 se
rect 5482 32761 5598 32773
tri 5598 32761 5610 32773 nw
tri 5732 32761 5744 32773 se
rect 5744 32761 14775 32773
rect 5482 32758 5595 32761
tri 5595 32758 5598 32761 nw
tri 5729 32758 5732 32761 se
rect 5732 32758 14775 32761
tri 5426 32717 5467 32758 se
rect 5467 32717 5554 32758
tri 5554 32717 5595 32758 nw
tri 5688 32717 5729 32758 se
rect 5729 32717 14775 32758
rect 14831 32717 14876 32773
rect 14932 32717 14977 32773
rect 15033 32717 15041 32773
tri 23431 32758 23451 32778 ne
rect 23451 32758 23501 32778
tri 23501 32758 23545 32802 sw
tri 23587 32758 23631 32802 ne
rect 23631 32770 23681 32802
tri 23681 32770 23713 32802 sw
tri 23767 32770 23799 32802 ne
rect 23799 32770 23861 32802
rect 23631 32762 23713 32770
tri 23713 32762 23721 32770 sw
tri 23799 32762 23807 32770 ne
rect 23807 32762 23861 32770
tri 23861 32762 23901 32802 sw
tri 23947 32762 23987 32802 ne
rect 23987 32776 24041 32802
tri 24041 32776 24067 32802 sw
tri 24127 32776 24153 32802 ne
rect 24153 32776 24221 32802
tri 24221 32776 24247 32802 sw
tri 24308 32776 24334 32802 ne
rect 24334 32776 24402 32802
tri 24402 32776 24428 32802 sw
rect 23987 32762 24067 32776
rect 23631 32758 23721 32762
tri 23721 32758 23725 32762 sw
tri 23807 32758 23811 32762 ne
rect 23811 32758 23901 32762
tri 23901 32758 23905 32762 sw
tri 23987 32758 23991 32762 ne
rect 23991 32758 24067 32762
tri 24067 32758 24085 32776 sw
tri 24153 32758 24171 32776 ne
rect 24171 32758 24247 32776
tri 24247 32758 24265 32776 sw
tri 24334 32758 24352 32776 ne
rect 24352 32758 24428 32776
tri 24428 32758 24446 32776 sw
tri 5406 32697 5426 32717 se
rect 5426 32697 5534 32717
tri 5534 32697 5554 32717 nw
tri 5683 32712 5688 32717 se
rect 5688 32712 15041 32717
rect 18133 32753 23365 32758
tri 5668 32697 5683 32712 se
rect 5683 32697 5819 32712
tri 5819 32697 5834 32712 nw
rect 18133 32697 18138 32753
rect 18194 32697 18218 32753
rect 18274 32748 23365 32753
tri 23365 32748 23375 32758 sw
tri 23451 32748 23461 32758 ne
rect 23461 32748 23545 32758
tri 23545 32748 23555 32758 sw
tri 23631 32748 23641 32758 ne
rect 23641 32748 23725 32758
tri 23725 32748 23735 32758 sw
tri 23811 32748 23821 32758 ne
rect 23821 32754 23905 32758
tri 23905 32754 23909 32758 sw
tri 23991 32754 23995 32758 ne
rect 23995 32754 24085 32758
rect 23821 32748 23909 32754
tri 23909 32748 23915 32754 sw
tri 23995 32748 24001 32754 ne
rect 24001 32748 24085 32754
tri 24085 32748 24095 32758 sw
tri 24171 32748 24181 32758 ne
rect 24181 32748 24265 32758
tri 24265 32748 24275 32758 sw
tri 24352 32748 24362 32758 ne
rect 24362 32748 24446 32758
tri 24446 32748 24456 32758 sw
rect 18274 32697 23375 32748
tri 5401 32692 5406 32697 se
rect 5406 32692 5529 32697
tri 5529 32692 5534 32697 nw
tri 5663 32692 5668 32697 se
rect 5668 32692 5814 32697
tri 5814 32692 5819 32697 nw
rect 18133 32694 23375 32697
tri 23375 32694 23429 32748 sw
tri 23461 32694 23515 32748 ne
rect 23515 32716 23555 32748
tri 23555 32716 23587 32748 sw
tri 23641 32716 23673 32748 ne
rect 23673 32716 23735 32748
rect 23515 32708 23587 32716
tri 23587 32708 23595 32716 sw
tri 23673 32708 23681 32716 ne
rect 23681 32708 23735 32716
tri 23735 32708 23775 32748 sw
tri 23821 32708 23861 32748 ne
rect 23861 32722 23915 32748
tri 23915 32722 23941 32748 sw
tri 24001 32722 24027 32748 ne
rect 24027 32722 24095 32748
tri 24095 32722 24121 32748 sw
tri 24181 32722 24207 32748 ne
rect 24207 32743 24275 32748
tri 24275 32743 24280 32748 sw
tri 24362 32743 24367 32748 ne
rect 24367 32743 24456 32748
rect 24207 32736 24280 32743
tri 24280 32736 24287 32743 sw
tri 24367 32736 24374 32743 ne
rect 24374 32736 24456 32743
tri 24456 32736 24468 32748 sw
rect 24207 32722 24287 32736
rect 23861 32708 23941 32722
tri 23941 32708 23955 32722 sw
tri 24027 32708 24041 32722 ne
rect 24041 32714 24121 32722
tri 24121 32714 24129 32722 sw
tri 24207 32714 24215 32722 ne
rect 24215 32714 24287 32722
rect 24041 32708 24129 32714
tri 24129 32708 24135 32714 sw
tri 24215 32708 24221 32714 ne
rect 24221 32708 24287 32714
tri 24287 32708 24315 32736 sw
tri 24374 32708 24402 32736 ne
rect 24402 32708 24468 32736
tri 24468 32708 24496 32736 sw
rect 23515 32694 23595 32708
tri 23595 32694 23609 32708 sw
tri 23681 32694 23695 32708 ne
rect 23695 32694 23775 32708
tri 23775 32694 23789 32708 sw
tri 23861 32694 23875 32708 ne
rect 23875 32694 23955 32708
tri 23955 32694 23969 32708 sw
tri 24041 32694 24055 32708 ne
rect 24055 32694 24135 32708
tri 24135 32694 24149 32708 sw
tri 24221 32694 24235 32708 ne
rect 24235 32694 24315 32708
tri 24315 32694 24329 32708 sw
tri 24402 32694 24416 32708 ne
rect 24416 32694 24496 32708
tri 24496 32694 24510 32708 sw
rect 18133 32692 23429 32694
tri 5375 32666 5401 32692 se
rect 5401 32666 5503 32692
tri 5503 32666 5529 32692 nw
tri 5637 32666 5663 32692 se
rect 5663 32666 5749 32692
rect 5375 32627 5464 32666
tri 5464 32627 5503 32666 nw
tri 5598 32627 5637 32666 se
rect 5637 32627 5749 32666
tri 5749 32627 5814 32692 nw
tri 23337 32627 23402 32692 ne
rect 23402 32662 23429 32692
tri 23429 32662 23461 32694 sw
tri 23515 32662 23547 32694 ne
rect 23547 32662 23609 32694
rect 23402 32654 23461 32662
tri 23461 32654 23469 32662 sw
tri 23547 32654 23555 32662 ne
rect 23555 32654 23609 32662
tri 23609 32654 23649 32694 sw
tri 23695 32654 23735 32694 ne
rect 23735 32676 23789 32694
tri 23789 32676 23807 32694 sw
tri 23875 32676 23893 32694 ne
rect 23893 32676 23969 32694
rect 23735 32668 23807 32676
tri 23807 32668 23815 32676 sw
tri 23893 32668 23901 32676 ne
rect 23901 32668 23969 32676
tri 23969 32668 23995 32694 sw
tri 24055 32668 24081 32694 ne
rect 24081 32682 24149 32694
tri 24149 32682 24161 32694 sw
tri 24235 32682 24247 32694 ne
rect 24247 32682 24329 32694
tri 24329 32682 24341 32694 sw
tri 24416 32682 24428 32694 ne
rect 24428 32682 24510 32694
tri 24510 32682 24522 32694 sw
rect 24081 32668 24161 32682
rect 23735 32654 23815 32668
tri 23815 32654 23829 32668 sw
tri 23901 32654 23915 32668 ne
rect 23915 32660 23995 32668
tri 23995 32660 24003 32668 sw
tri 24081 32660 24089 32668 ne
rect 24089 32660 24161 32668
rect 23915 32654 24003 32660
tri 24003 32654 24009 32660 sw
tri 24089 32654 24095 32660 ne
rect 24095 32654 24161 32660
tri 24161 32654 24189 32682 sw
tri 24247 32654 24275 32682 ne
rect 24275 32654 24341 32682
tri 24341 32654 24369 32682 sw
tri 24428 32654 24456 32682 ne
rect 24456 32654 24522 32682
tri 24522 32654 24550 32682 sw
rect 23402 32627 23469 32654
tri 5334 29432 5375 29473 se
rect 5375 29432 5441 32627
tri 5441 32604 5464 32627 nw
tri 5575 32604 5598 32627 se
rect 5598 32604 5722 32627
tri 5571 32600 5575 32604 se
rect 5575 32600 5722 32604
tri 5722 32600 5749 32627 nw
tri 23402 32600 23429 32627 ne
rect 23429 32600 23469 32627
tri 23469 32600 23523 32654 sw
tri 23555 32600 23609 32654 ne
rect 23609 32622 23649 32654
tri 23649 32622 23681 32654 sw
tri 23735 32622 23767 32654 ne
rect 23767 32622 23829 32654
rect 23609 32614 23681 32622
tri 23681 32614 23689 32622 sw
tri 23767 32614 23775 32622 ne
rect 23775 32614 23829 32622
tri 23829 32614 23869 32654 sw
tri 23915 32614 23955 32654 ne
rect 23955 32628 24009 32654
tri 24009 32628 24035 32654 sw
tri 24095 32628 24121 32654 ne
rect 24121 32628 24189 32654
tri 24189 32628 24215 32654 sw
tri 24275 32628 24301 32654 ne
rect 24301 32649 24369 32654
tri 24369 32649 24374 32654 sw
tri 24456 32649 24461 32654 ne
rect 24461 32649 24550 32654
rect 24301 32642 24374 32649
tri 24374 32642 24381 32649 sw
tri 24461 32642 24468 32649 ne
rect 24468 32642 24550 32649
tri 24550 32642 24562 32654 sw
rect 24301 32628 24381 32642
rect 23955 32614 24035 32628
tri 24035 32614 24049 32628 sw
tri 24121 32614 24135 32628 ne
rect 24135 32620 24215 32628
tri 24215 32620 24223 32628 sw
tri 24301 32620 24309 32628 ne
rect 24309 32620 24381 32628
rect 24135 32614 24223 32620
tri 24223 32614 24229 32620 sw
tri 24309 32614 24315 32620 ne
rect 24315 32614 24381 32620
tri 24381 32614 24409 32642 sw
tri 24468 32614 24496 32642 ne
rect 24496 32614 24562 32642
tri 24562 32614 24590 32642 sw
rect 23609 32600 23689 32614
tri 23689 32600 23703 32614 sw
tri 23775 32600 23789 32614 ne
rect 23789 32600 23869 32614
tri 23869 32600 23883 32614 sw
tri 23955 32600 23969 32614 ne
rect 23969 32600 24049 32614
tri 24049 32600 24063 32614 sw
tri 24135 32600 24149 32614 ne
rect 24149 32600 24229 32614
tri 24229 32600 24243 32614 sw
tri 24315 32600 24329 32614 ne
rect 24329 32600 24409 32614
tri 24409 32600 24423 32614 sw
tri 24496 32600 24510 32614 ne
rect 24510 32600 24590 32614
tri 24590 32600 24604 32614 sw
tri 5295 29393 5334 29432 se
rect 5334 29393 5441 29432
tri 5501 32530 5571 32600 se
rect 5571 32530 5652 32600
tri 5652 32530 5722 32600 nw
tri 23429 32530 23499 32600 ne
rect 23499 32568 23523 32600
tri 23523 32568 23555 32600 sw
tri 23609 32568 23641 32600 ne
rect 23641 32568 23703 32600
rect 23499 32560 23555 32568
tri 23555 32560 23563 32568 sw
tri 23641 32560 23649 32568 ne
rect 23649 32560 23703 32568
tri 23703 32560 23743 32600 sw
tri 23789 32560 23829 32600 ne
rect 23829 32582 23883 32600
tri 23883 32582 23901 32600 sw
tri 23969 32582 23987 32600 ne
rect 23987 32582 24063 32600
rect 23829 32574 23901 32582
tri 23901 32574 23909 32582 sw
tri 23987 32574 23995 32582 ne
rect 23995 32574 24063 32582
tri 24063 32574 24089 32600 sw
tri 24149 32574 24175 32600 ne
rect 24175 32588 24243 32600
tri 24243 32588 24255 32600 sw
tri 24329 32588 24341 32600 ne
rect 24341 32588 24423 32600
tri 24423 32588 24435 32600 sw
tri 24510 32588 24522 32600 ne
rect 24522 32588 24604 32600
tri 24604 32588 24616 32600 sw
rect 24175 32574 24255 32588
rect 23829 32560 23909 32574
tri 23909 32560 23923 32574 sw
tri 23995 32560 24009 32574 ne
rect 24009 32566 24089 32574
tri 24089 32566 24097 32574 sw
tri 24175 32566 24183 32574 ne
rect 24183 32566 24255 32574
rect 24009 32560 24097 32566
tri 24097 32560 24103 32566 sw
tri 24183 32560 24189 32566 ne
rect 24189 32560 24255 32566
tri 24255 32560 24283 32588 sw
tri 24341 32560 24369 32588 ne
rect 24369 32560 24435 32588
tri 24435 32560 24463 32588 sw
tri 24522 32560 24550 32588 ne
rect 24550 32560 24616 32588
tri 24616 32560 24644 32588 sw
rect 23499 32530 23563 32560
rect 5501 32506 5628 32530
tri 5628 32506 5652 32530 nw
tri 23499 32506 23523 32530 ne
rect 23523 32506 23563 32530
tri 23563 32506 23617 32560 sw
tri 23649 32506 23703 32560 ne
rect 23703 32528 23743 32560
tri 23743 32528 23775 32560 sw
tri 23829 32528 23861 32560 ne
rect 23861 32528 23923 32560
rect 23703 32520 23775 32528
tri 23775 32520 23783 32528 sw
tri 23861 32520 23869 32528 ne
rect 23869 32520 23923 32528
tri 23923 32520 23963 32560 sw
tri 24009 32520 24049 32560 ne
rect 24049 32534 24103 32560
tri 24103 32534 24129 32560 sw
tri 24189 32534 24215 32560 ne
rect 24215 32534 24283 32560
tri 24283 32534 24309 32560 sw
tri 24369 32534 24395 32560 ne
rect 24395 32555 24463 32560
tri 24463 32555 24468 32560 sw
tri 24550 32555 24555 32560 ne
rect 24555 32555 24644 32560
rect 24395 32548 24468 32555
tri 24468 32548 24475 32555 sw
tri 24555 32548 24562 32555 ne
rect 24562 32548 24644 32555
tri 24644 32548 24656 32560 sw
rect 24395 32534 24475 32548
rect 24049 32520 24129 32534
tri 24129 32520 24143 32534 sw
tri 24215 32520 24229 32534 ne
rect 24229 32526 24309 32534
tri 24309 32526 24317 32534 sw
tri 24395 32526 24403 32534 ne
rect 24403 32526 24475 32534
rect 24229 32520 24317 32526
tri 24317 32520 24323 32526 sw
tri 24403 32520 24409 32526 ne
rect 24409 32520 24475 32526
tri 24475 32520 24503 32548 sw
tri 24562 32520 24590 32548 ne
rect 24590 32520 24656 32548
tri 24656 32520 24684 32548 sw
rect 23703 32506 23783 32520
tri 23783 32506 23797 32520 sw
tri 23869 32506 23883 32520 ne
rect 23883 32506 23963 32520
tri 23963 32506 23977 32520 sw
tri 24049 32506 24063 32520 ne
rect 24063 32506 24143 32520
tri 24143 32506 24157 32520 sw
tri 24229 32506 24243 32520 ne
rect 24243 32506 24323 32520
tri 24323 32506 24337 32520 sw
tri 24409 32506 24423 32520 ne
rect 24423 32506 24503 32520
tri 24503 32506 24517 32520 sw
tri 24590 32506 24604 32520 ne
rect 24604 32506 24684 32520
tri 24684 32506 24698 32520 sw
rect 5501 29493 5567 32506
tri 5567 32445 5628 32506 nw
tri 23523 32445 23584 32506 ne
rect 23584 32474 23617 32506
tri 23617 32474 23649 32506 sw
tri 23703 32474 23735 32506 ne
rect 23735 32474 23797 32506
rect 23584 32466 23649 32474
tri 23649 32466 23657 32474 sw
tri 23735 32466 23743 32474 ne
rect 23743 32466 23797 32474
tri 23797 32466 23837 32506 sw
tri 23883 32466 23923 32506 ne
rect 23923 32488 23977 32506
tri 23977 32488 23995 32506 sw
tri 24063 32488 24081 32506 ne
rect 24081 32488 24157 32506
rect 23923 32480 23995 32488
tri 23995 32480 24003 32488 sw
tri 24081 32480 24089 32488 ne
rect 24089 32480 24157 32488
tri 24157 32480 24183 32506 sw
tri 24243 32480 24269 32506 ne
rect 24269 32494 24337 32506
tri 24337 32494 24349 32506 sw
tri 24423 32494 24435 32506 ne
rect 24435 32494 24517 32506
tri 24517 32494 24529 32506 sw
tri 24604 32494 24616 32506 ne
rect 24616 32494 24698 32506
tri 24698 32494 24710 32506 sw
rect 24269 32480 24349 32494
rect 23923 32466 24003 32480
tri 24003 32466 24017 32480 sw
tri 24089 32466 24103 32480 ne
rect 24103 32472 24183 32480
tri 24183 32472 24191 32480 sw
tri 24269 32472 24277 32480 ne
rect 24277 32472 24349 32480
rect 24103 32466 24191 32472
tri 24191 32466 24197 32472 sw
tri 24277 32466 24283 32472 ne
rect 24283 32466 24349 32472
tri 24349 32466 24377 32494 sw
tri 24435 32466 24463 32494 ne
rect 24463 32466 24529 32494
tri 24529 32466 24557 32494 sw
tri 24616 32466 24644 32494 ne
rect 24644 32466 24710 32494
tri 24710 32466 24738 32494 sw
rect 23584 32445 23657 32466
tri 23584 32412 23617 32445 ne
rect 23617 32412 23657 32445
tri 23657 32412 23711 32466 sw
tri 23743 32412 23797 32466 ne
rect 23797 32434 23837 32466
tri 23837 32434 23869 32466 sw
tri 23923 32434 23955 32466 ne
rect 23955 32434 24017 32466
rect 23797 32426 23869 32434
tri 23869 32426 23877 32434 sw
tri 23955 32426 23963 32434 ne
rect 23963 32426 24017 32434
tri 24017 32426 24057 32466 sw
tri 24103 32426 24143 32466 ne
rect 24143 32440 24197 32466
tri 24197 32440 24223 32466 sw
tri 24283 32440 24309 32466 ne
rect 24309 32440 24377 32466
tri 24377 32440 24403 32466 sw
tri 24463 32440 24489 32466 ne
rect 24489 32461 24557 32466
tri 24557 32461 24562 32466 sw
tri 24644 32461 24649 32466 ne
rect 24649 32461 24738 32466
rect 24489 32454 24562 32461
tri 24562 32454 24569 32461 sw
tri 24649 32454 24656 32461 ne
rect 24656 32454 24738 32461
tri 24738 32454 24750 32466 sw
rect 24489 32440 24569 32454
rect 24143 32426 24223 32440
tri 24223 32426 24237 32440 sw
tri 24309 32426 24323 32440 ne
rect 24323 32432 24403 32440
tri 24403 32432 24411 32440 sw
tri 24489 32432 24497 32440 ne
rect 24497 32432 24569 32440
rect 24323 32426 24411 32432
tri 24411 32426 24417 32432 sw
tri 24497 32426 24503 32432 ne
rect 24503 32426 24569 32432
tri 24569 32426 24597 32454 sw
tri 24656 32426 24684 32454 ne
rect 24684 32426 24750 32454
tri 24750 32426 24778 32454 sw
rect 23797 32412 23877 32426
tri 23877 32412 23891 32426 sw
tri 23963 32412 23977 32426 ne
rect 23977 32412 24057 32426
tri 24057 32412 24071 32426 sw
tri 24143 32412 24157 32426 ne
rect 24157 32412 24237 32426
tri 24237 32412 24251 32426 sw
tri 24323 32412 24337 32426 ne
rect 24337 32412 24417 32426
tri 24417 32412 24431 32426 sw
tri 24503 32412 24517 32426 ne
rect 24517 32412 24597 32426
tri 24597 32412 24611 32426 sw
tri 24684 32412 24698 32426 ne
rect 24698 32412 24778 32426
tri 24778 32412 24792 32426 sw
tri 23617 32318 23711 32412 ne
tri 23711 32380 23743 32412 sw
tri 23797 32380 23829 32412 ne
rect 23829 32380 23891 32412
rect 23711 32372 23743 32380
tri 23743 32372 23751 32380 sw
tri 23829 32372 23837 32380 ne
rect 23837 32372 23891 32380
tri 23891 32372 23931 32412 sw
tri 23977 32372 24017 32412 ne
rect 24017 32394 24071 32412
tri 24071 32394 24089 32412 sw
tri 24157 32394 24175 32412 ne
rect 24175 32394 24251 32412
rect 24017 32386 24089 32394
tri 24089 32386 24097 32394 sw
tri 24175 32386 24183 32394 ne
rect 24183 32386 24251 32394
tri 24251 32386 24277 32412 sw
tri 24337 32386 24363 32412 ne
rect 24363 32400 24431 32412
tri 24431 32400 24443 32412 sw
tri 24517 32400 24529 32412 ne
rect 24529 32400 24611 32412
tri 24611 32400 24623 32412 sw
tri 24698 32400 24710 32412 ne
rect 24710 32400 24792 32412
tri 24792 32400 24804 32412 sw
rect 24363 32386 24443 32400
rect 24017 32372 24097 32386
tri 24097 32372 24111 32386 sw
tri 24183 32372 24197 32386 ne
rect 24197 32378 24277 32386
tri 24277 32378 24285 32386 sw
tri 24363 32378 24371 32386 ne
rect 24371 32378 24443 32386
rect 24197 32372 24285 32378
tri 24285 32372 24291 32378 sw
tri 24371 32372 24377 32378 ne
rect 24377 32372 24443 32378
tri 24443 32372 24471 32400 sw
tri 24529 32372 24557 32400 ne
rect 24557 32372 24623 32400
tri 24623 32372 24651 32400 sw
tri 24710 32372 24738 32400 ne
rect 24738 32372 24804 32400
tri 24804 32372 24832 32400 sw
rect 23711 32318 23751 32372
tri 23751 32318 23805 32372 sw
tri 23837 32318 23891 32372 ne
rect 23891 32340 23931 32372
tri 23931 32340 23963 32372 sw
tri 24017 32340 24049 32372 ne
rect 24049 32340 24111 32372
rect 23891 32332 23963 32340
tri 23963 32332 23971 32340 sw
tri 24049 32332 24057 32340 ne
rect 24057 32332 24111 32340
tri 24111 32332 24151 32372 sw
tri 24197 32332 24237 32372 ne
rect 24237 32346 24291 32372
tri 24291 32346 24317 32372 sw
tri 24377 32346 24403 32372 ne
rect 24403 32346 24471 32372
tri 24471 32346 24497 32372 sw
tri 24557 32346 24583 32372 ne
rect 24583 32367 24651 32372
tri 24651 32367 24656 32372 sw
tri 24738 32367 24743 32372 ne
rect 24743 32367 24832 32372
rect 24583 32360 24656 32367
tri 24656 32360 24663 32367 sw
tri 24743 32360 24750 32367 ne
rect 24750 32360 24832 32367
tri 24832 32360 24844 32372 sw
rect 24583 32346 24663 32360
rect 24237 32332 24317 32346
tri 24317 32332 24331 32346 sw
tri 24403 32332 24417 32346 ne
rect 24417 32338 24497 32346
tri 24497 32338 24505 32346 sw
tri 24583 32338 24591 32346 ne
rect 24591 32338 24663 32346
rect 24417 32332 24505 32338
tri 24505 32332 24511 32338 sw
tri 24591 32332 24597 32338 ne
rect 24597 32332 24663 32338
tri 24663 32332 24691 32360 sw
tri 24750 32332 24778 32360 ne
rect 24778 32332 24844 32360
tri 24844 32332 24872 32360 sw
rect 23891 32318 23971 32332
tri 23971 32318 23985 32332 sw
tri 24057 32318 24071 32332 ne
rect 24071 32318 24151 32332
tri 24151 32318 24165 32332 sw
tri 24237 32318 24251 32332 ne
rect 24251 32318 24331 32332
tri 24331 32318 24345 32332 sw
tri 24417 32318 24431 32332 ne
rect 24431 32318 24511 32332
tri 24511 32318 24525 32332 sw
tri 24597 32318 24611 32332 ne
rect 24611 32318 24691 32332
tri 24691 32318 24705 32332 sw
tri 24778 32318 24792 32332 ne
rect 24792 32318 24872 32332
tri 24872 32318 24886 32332 sw
tri 23711 32224 23805 32318 ne
tri 23805 32286 23837 32318 sw
tri 23891 32286 23923 32318 ne
rect 23923 32286 23985 32318
rect 23805 32278 23837 32286
tri 23837 32278 23845 32286 sw
tri 23923 32278 23931 32286 ne
rect 23931 32278 23985 32286
tri 23985 32278 24025 32318 sw
tri 24071 32278 24111 32318 ne
rect 24111 32300 24165 32318
tri 24165 32300 24183 32318 sw
tri 24251 32300 24269 32318 ne
rect 24269 32300 24345 32318
rect 24111 32292 24183 32300
tri 24183 32292 24191 32300 sw
tri 24269 32292 24277 32300 ne
rect 24277 32292 24345 32300
tri 24345 32292 24371 32318 sw
tri 24431 32292 24457 32318 ne
rect 24457 32306 24525 32318
tri 24525 32306 24537 32318 sw
tri 24611 32306 24623 32318 ne
rect 24623 32306 24705 32318
tri 24705 32306 24717 32318 sw
tri 24792 32306 24804 32318 ne
rect 24804 32306 24886 32318
tri 24886 32306 24898 32318 sw
rect 24457 32292 24537 32306
rect 24111 32278 24191 32292
tri 24191 32278 24205 32292 sw
tri 24277 32278 24291 32292 ne
rect 24291 32284 24371 32292
tri 24371 32284 24379 32292 sw
tri 24457 32284 24465 32292 ne
rect 24465 32284 24537 32292
rect 24291 32278 24379 32284
tri 24379 32278 24385 32284 sw
tri 24465 32278 24471 32284 ne
rect 24471 32278 24537 32284
tri 24537 32278 24565 32306 sw
tri 24623 32278 24651 32306 ne
rect 24651 32278 24717 32306
tri 24717 32278 24745 32306 sw
tri 24804 32278 24832 32306 ne
rect 24832 32278 24898 32306
tri 24898 32278 24926 32306 sw
rect 23805 32224 23845 32278
tri 23845 32224 23899 32278 sw
tri 23931 32224 23985 32278 ne
rect 23985 32246 24025 32278
tri 24025 32246 24057 32278 sw
tri 24111 32246 24143 32278 ne
rect 24143 32246 24205 32278
rect 23985 32238 24057 32246
tri 24057 32238 24065 32246 sw
tri 24143 32238 24151 32246 ne
rect 24151 32238 24205 32246
tri 24205 32238 24245 32278 sw
tri 24291 32238 24331 32278 ne
rect 24331 32252 24385 32278
tri 24385 32252 24411 32278 sw
tri 24471 32252 24497 32278 ne
rect 24497 32252 24565 32278
tri 24565 32252 24591 32278 sw
tri 24651 32252 24677 32278 ne
rect 24677 32273 24745 32278
tri 24745 32273 24750 32278 sw
tri 24832 32273 24837 32278 ne
rect 24837 32273 24926 32278
rect 24677 32266 24750 32273
tri 24750 32266 24757 32273 sw
tri 24837 32266 24844 32273 ne
rect 24844 32266 24926 32273
tri 24926 32266 24938 32278 sw
rect 24677 32252 24757 32266
rect 24331 32238 24411 32252
tri 24411 32238 24425 32252 sw
tri 24497 32238 24511 32252 ne
rect 24511 32244 24591 32252
tri 24591 32244 24599 32252 sw
tri 24677 32244 24685 32252 ne
rect 24685 32244 24757 32252
rect 24511 32238 24599 32244
tri 24599 32238 24605 32244 sw
tri 24685 32238 24691 32244 ne
rect 24691 32238 24757 32244
tri 24757 32238 24785 32266 sw
tri 24844 32238 24872 32266 ne
rect 24872 32238 24938 32266
tri 24938 32238 24966 32266 sw
rect 23985 32224 24065 32238
tri 24065 32224 24079 32238 sw
tri 24151 32224 24165 32238 ne
rect 24165 32224 24245 32238
tri 24245 32224 24259 32238 sw
tri 24331 32224 24345 32238 ne
rect 24345 32224 24425 32238
tri 24425 32224 24439 32238 sw
tri 24511 32224 24525 32238 ne
rect 24525 32224 24605 32238
tri 24605 32224 24619 32238 sw
tri 24691 32224 24705 32238 ne
rect 24705 32224 24785 32238
tri 24785 32224 24799 32238 sw
tri 24872 32224 24886 32238 ne
rect 24886 32224 24966 32238
tri 24966 32224 24980 32238 sw
tri 23805 32130 23899 32224 ne
tri 23899 32192 23931 32224 sw
tri 23985 32192 24017 32224 ne
rect 24017 32192 24079 32224
rect 23899 32184 23931 32192
tri 23931 32184 23939 32192 sw
tri 24017 32184 24025 32192 ne
rect 24025 32184 24079 32192
tri 24079 32184 24119 32224 sw
tri 24165 32184 24205 32224 ne
rect 24205 32206 24259 32224
tri 24259 32206 24277 32224 sw
tri 24345 32206 24363 32224 ne
rect 24363 32206 24439 32224
rect 24205 32198 24277 32206
tri 24277 32198 24285 32206 sw
tri 24363 32198 24371 32206 ne
rect 24371 32198 24439 32206
tri 24439 32198 24465 32224 sw
tri 24525 32198 24551 32224 ne
rect 24551 32212 24619 32224
tri 24619 32212 24631 32224 sw
tri 24705 32212 24717 32224 ne
rect 24717 32212 24799 32224
tri 24799 32212 24811 32224 sw
tri 24886 32212 24898 32224 ne
rect 24898 32212 24980 32224
tri 24980 32212 24992 32224 sw
rect 24551 32198 24631 32212
rect 24205 32184 24285 32198
tri 24285 32184 24299 32198 sw
tri 24371 32184 24385 32198 ne
rect 24385 32190 24465 32198
tri 24465 32190 24473 32198 sw
tri 24551 32190 24559 32198 ne
rect 24559 32190 24631 32198
rect 24385 32184 24473 32190
tri 24473 32184 24479 32190 sw
tri 24559 32184 24565 32190 ne
rect 24565 32184 24631 32190
tri 24631 32184 24659 32212 sw
tri 24717 32184 24745 32212 ne
rect 24745 32184 24811 32212
tri 24811 32184 24839 32212 sw
tri 24898 32184 24926 32212 ne
rect 24926 32184 24992 32212
tri 24992 32184 25020 32212 sw
rect 23899 32130 23939 32184
tri 23939 32130 23993 32184 sw
tri 24025 32130 24079 32184 ne
rect 24079 32152 24119 32184
tri 24119 32152 24151 32184 sw
tri 24205 32152 24237 32184 ne
rect 24237 32152 24299 32184
rect 24079 32144 24151 32152
tri 24151 32144 24159 32152 sw
tri 24237 32144 24245 32152 ne
rect 24245 32144 24299 32152
tri 24299 32144 24339 32184 sw
tri 24385 32144 24425 32184 ne
rect 24425 32158 24479 32184
tri 24479 32158 24505 32184 sw
tri 24565 32158 24591 32184 ne
rect 24591 32158 24659 32184
tri 24659 32158 24685 32184 sw
tri 24745 32158 24771 32184 ne
rect 24771 32179 24839 32184
tri 24839 32179 24844 32184 sw
tri 24926 32179 24931 32184 ne
rect 24931 32179 25020 32184
rect 24771 32172 24844 32179
tri 24844 32172 24851 32179 sw
tri 24931 32172 24938 32179 ne
rect 24938 32172 25020 32179
tri 25020 32172 25032 32184 sw
rect 24771 32158 24851 32172
rect 24425 32144 24505 32158
tri 24505 32144 24519 32158 sw
tri 24591 32144 24605 32158 ne
rect 24605 32150 24685 32158
tri 24685 32150 24693 32158 sw
tri 24771 32150 24779 32158 ne
rect 24779 32150 24851 32158
rect 24605 32144 24693 32150
tri 24693 32144 24699 32150 sw
tri 24779 32144 24785 32150 ne
rect 24785 32144 24851 32150
tri 24851 32144 24879 32172 sw
tri 24938 32144 24966 32172 ne
rect 24966 32144 25032 32172
tri 25032 32144 25060 32172 sw
rect 24079 32130 24159 32144
tri 24159 32130 24173 32144 sw
tri 24245 32130 24259 32144 ne
rect 24259 32130 24339 32144
tri 24339 32130 24353 32144 sw
tri 24425 32130 24439 32144 ne
rect 24439 32130 24519 32144
tri 24519 32130 24533 32144 sw
tri 24605 32130 24619 32144 ne
rect 24619 32130 24699 32144
tri 24699 32130 24713 32144 sw
tri 24785 32130 24799 32144 ne
rect 24799 32130 24879 32144
tri 24879 32130 24893 32144 sw
tri 24966 32130 24980 32144 ne
rect 24980 32130 25060 32144
tri 25060 32130 25074 32144 sw
tri 23899 32036 23993 32130 ne
tri 23993 32098 24025 32130 sw
tri 24079 32098 24111 32130 ne
rect 24111 32098 24173 32130
rect 23993 32090 24025 32098
tri 24025 32090 24033 32098 sw
tri 24111 32090 24119 32098 ne
rect 24119 32090 24173 32098
tri 24173 32090 24213 32130 sw
tri 24259 32090 24299 32130 ne
rect 24299 32112 24353 32130
tri 24353 32112 24371 32130 sw
tri 24439 32112 24457 32130 ne
rect 24457 32112 24533 32130
rect 24299 32104 24371 32112
tri 24371 32104 24379 32112 sw
tri 24457 32104 24465 32112 ne
rect 24465 32104 24533 32112
tri 24533 32104 24559 32130 sw
tri 24619 32104 24645 32130 ne
rect 24645 32118 24713 32130
tri 24713 32118 24725 32130 sw
tri 24799 32118 24811 32130 ne
rect 24811 32118 24893 32130
tri 24893 32118 24905 32130 sw
tri 24980 32118 24992 32130 ne
rect 24992 32118 25074 32130
tri 25074 32118 25086 32130 sw
rect 24645 32104 24725 32118
rect 24299 32090 24379 32104
tri 24379 32090 24393 32104 sw
tri 24465 32090 24479 32104 ne
rect 24479 32096 24559 32104
tri 24559 32096 24567 32104 sw
tri 24645 32096 24653 32104 ne
rect 24653 32096 24725 32104
rect 24479 32090 24567 32096
tri 24567 32090 24573 32096 sw
tri 24653 32090 24659 32096 ne
rect 24659 32090 24725 32096
tri 24725 32090 24753 32118 sw
tri 24811 32090 24839 32118 ne
rect 24839 32090 24905 32118
tri 24905 32090 24933 32118 sw
tri 24992 32090 25020 32118 ne
rect 25020 32090 25086 32118
tri 25086 32090 25114 32118 sw
rect 23993 32036 24033 32090
tri 24033 32036 24087 32090 sw
tri 24119 32036 24173 32090 ne
rect 24173 32058 24213 32090
tri 24213 32058 24245 32090 sw
tri 24299 32058 24331 32090 ne
rect 24331 32058 24393 32090
rect 24173 32050 24245 32058
tri 24245 32050 24253 32058 sw
tri 24331 32050 24339 32058 ne
rect 24339 32050 24393 32058
tri 24393 32050 24433 32090 sw
tri 24479 32050 24519 32090 ne
rect 24519 32064 24573 32090
tri 24573 32064 24599 32090 sw
tri 24659 32064 24685 32090 ne
rect 24685 32064 24753 32090
tri 24753 32064 24779 32090 sw
tri 24839 32064 24865 32090 ne
rect 24865 32085 24933 32090
tri 24933 32085 24938 32090 sw
tri 25020 32085 25025 32090 ne
rect 25025 32085 25114 32090
rect 24865 32078 24938 32085
tri 24938 32078 24945 32085 sw
tri 25025 32078 25032 32085 ne
rect 25032 32078 25114 32085
tri 25114 32078 25126 32090 sw
rect 24865 32064 24945 32078
rect 24519 32050 24599 32064
tri 24599 32050 24613 32064 sw
tri 24685 32050 24699 32064 ne
rect 24699 32056 24779 32064
tri 24779 32056 24787 32064 sw
tri 24865 32056 24873 32064 ne
rect 24873 32056 24945 32064
rect 24699 32050 24787 32056
tri 24787 32050 24793 32056 sw
tri 24873 32050 24879 32056 ne
rect 24879 32050 24945 32056
tri 24945 32050 24973 32078 sw
tri 25032 32050 25060 32078 ne
rect 25060 32050 25126 32078
tri 25126 32050 25154 32078 sw
rect 24173 32036 24253 32050
tri 24253 32036 24267 32050 sw
tri 24339 32036 24353 32050 ne
rect 24353 32036 24433 32050
tri 24433 32036 24447 32050 sw
tri 24519 32036 24533 32050 ne
rect 24533 32036 24613 32050
tri 24613 32036 24627 32050 sw
tri 24699 32036 24713 32050 ne
rect 24713 32036 24793 32050
tri 24793 32036 24807 32050 sw
tri 24879 32036 24893 32050 ne
rect 24893 32036 24973 32050
tri 24973 32036 24987 32050 sw
tri 25060 32036 25074 32050 ne
rect 25074 32036 25154 32050
tri 25154 32036 25168 32050 sw
tri 23993 31942 24087 32036 ne
tri 24087 32004 24119 32036 sw
tri 24173 32004 24205 32036 ne
rect 24205 32004 24267 32036
rect 24087 31996 24119 32004
tri 24119 31996 24127 32004 sw
tri 24205 31996 24213 32004 ne
rect 24213 31996 24267 32004
tri 24267 31996 24307 32036 sw
tri 24353 31996 24393 32036 ne
rect 24393 32018 24447 32036
tri 24447 32018 24465 32036 sw
tri 24533 32018 24551 32036 ne
rect 24551 32018 24627 32036
rect 24393 32010 24465 32018
tri 24465 32010 24473 32018 sw
tri 24551 32010 24559 32018 ne
rect 24559 32010 24627 32018
tri 24627 32010 24653 32036 sw
tri 24713 32010 24739 32036 ne
rect 24739 32024 24807 32036
tri 24807 32024 24819 32036 sw
tri 24893 32024 24905 32036 ne
rect 24905 32024 24987 32036
tri 24987 32024 24999 32036 sw
tri 25074 32024 25086 32036 ne
rect 25086 32024 25168 32036
tri 25168 32024 25180 32036 sw
rect 24739 32010 24819 32024
rect 24393 31996 24473 32010
tri 24473 31996 24487 32010 sw
tri 24559 31996 24573 32010 ne
rect 24573 32002 24653 32010
tri 24653 32002 24661 32010 sw
tri 24739 32002 24747 32010 ne
rect 24747 32002 24819 32010
rect 24573 31996 24661 32002
tri 24661 31996 24667 32002 sw
tri 24747 31996 24753 32002 ne
rect 24753 31996 24819 32002
tri 24819 31996 24847 32024 sw
tri 24905 31996 24933 32024 ne
rect 24933 31996 24999 32024
tri 24999 31996 25027 32024 sw
tri 25086 31996 25114 32024 ne
rect 25114 31996 25180 32024
tri 25180 31996 25208 32024 sw
rect 24087 31942 24127 31996
tri 24127 31942 24181 31996 sw
tri 24213 31942 24267 31996 ne
rect 24267 31964 24307 31996
tri 24307 31964 24339 31996 sw
tri 24393 31964 24425 31996 ne
rect 24425 31964 24487 31996
rect 24267 31956 24339 31964
tri 24339 31956 24347 31964 sw
tri 24425 31956 24433 31964 ne
rect 24433 31956 24487 31964
tri 24487 31956 24527 31996 sw
tri 24573 31956 24613 31996 ne
rect 24613 31970 24667 31996
tri 24667 31970 24693 31996 sw
tri 24753 31970 24779 31996 ne
rect 24779 31970 24847 31996
tri 24847 31970 24873 31996 sw
tri 24933 31970 24959 31996 ne
rect 24959 31991 25027 31996
tri 25027 31991 25032 31996 sw
tri 25114 31991 25119 31996 ne
rect 25119 31991 25208 31996
rect 24959 31984 25032 31991
tri 25032 31984 25039 31991 sw
tri 25119 31984 25126 31991 ne
rect 25126 31984 25208 31991
tri 25208 31984 25220 31996 sw
rect 24959 31970 25039 31984
rect 24613 31956 24693 31970
tri 24693 31956 24707 31970 sw
tri 24779 31956 24793 31970 ne
rect 24793 31962 24873 31970
tri 24873 31962 24881 31970 sw
tri 24959 31962 24967 31970 ne
rect 24967 31962 25039 31970
rect 24793 31956 24881 31962
tri 24881 31956 24887 31962 sw
tri 24967 31956 24973 31962 ne
rect 24973 31956 25039 31962
tri 25039 31956 25067 31984 sw
tri 25126 31956 25154 31984 ne
rect 24267 31942 24347 31956
tri 24347 31942 24361 31956 sw
tri 24433 31942 24447 31956 ne
rect 24447 31942 24527 31956
tri 24527 31942 24541 31956 sw
tri 24613 31942 24627 31956 ne
rect 24627 31942 24707 31956
tri 24707 31942 24721 31956 sw
tri 24793 31942 24807 31956 ne
rect 24807 31942 24887 31956
tri 24887 31942 24901 31956 sw
tri 24973 31942 24987 31956 ne
rect 24987 31942 25067 31956
tri 25067 31942 25081 31956 sw
tri 24087 31848 24181 31942 ne
tri 24181 31910 24213 31942 sw
tri 24267 31910 24299 31942 ne
rect 24299 31910 24361 31942
rect 24181 31902 24213 31910
tri 24213 31902 24221 31910 sw
tri 24299 31902 24307 31910 ne
rect 24307 31902 24361 31910
tri 24361 31902 24401 31942 sw
tri 24447 31902 24487 31942 ne
rect 24487 31924 24541 31942
tri 24541 31924 24559 31942 sw
tri 24627 31924 24645 31942 ne
rect 24645 31924 24721 31942
rect 24487 31916 24559 31924
tri 24559 31916 24567 31924 sw
tri 24645 31916 24653 31924 ne
rect 24653 31916 24721 31924
tri 24721 31916 24747 31942 sw
tri 24807 31916 24833 31942 ne
rect 24833 31930 24901 31942
tri 24901 31930 24913 31942 sw
tri 24987 31930 24999 31942 ne
rect 24999 31930 25081 31942
tri 25081 31930 25093 31942 sw
rect 24833 31916 24913 31930
rect 24487 31902 24567 31916
tri 24567 31902 24581 31916 sw
tri 24653 31902 24667 31916 ne
rect 24667 31908 24747 31916
tri 24747 31908 24755 31916 sw
tri 24833 31908 24841 31916 ne
rect 24841 31908 24913 31916
rect 24667 31902 24755 31908
tri 24755 31902 24761 31908 sw
tri 24841 31902 24847 31908 ne
rect 24847 31902 24913 31908
tri 24913 31902 24941 31930 sw
tri 24999 31902 25027 31930 ne
rect 24181 31848 24221 31902
tri 24221 31848 24275 31902 sw
tri 24307 31848 24361 31902 ne
rect 24361 31870 24401 31902
tri 24401 31870 24433 31902 sw
tri 24487 31870 24519 31902 ne
rect 24519 31870 24581 31902
rect 24361 31862 24433 31870
tri 24433 31862 24441 31870 sw
tri 24519 31862 24527 31870 ne
rect 24527 31862 24581 31870
tri 24581 31862 24621 31902 sw
tri 24667 31862 24707 31902 ne
rect 24707 31876 24761 31902
tri 24761 31876 24787 31902 sw
tri 24847 31876 24873 31902 ne
rect 24873 31876 24941 31902
tri 24941 31876 24967 31902 sw
rect 24707 31862 24787 31876
tri 24787 31862 24801 31876 sw
tri 24873 31862 24887 31876 ne
rect 24887 31862 24967 31876
rect 24361 31848 24441 31862
tri 24441 31848 24455 31862 sw
tri 24527 31848 24541 31862 ne
rect 24541 31848 24621 31862
tri 24621 31848 24635 31862 sw
tri 24707 31848 24721 31862 ne
rect 24721 31848 24801 31862
tri 24801 31848 24815 31862 sw
tri 24887 31848 24901 31862 ne
tri 24181 31754 24275 31848 ne
tri 24275 31816 24307 31848 sw
tri 24361 31816 24393 31848 ne
rect 24393 31816 24455 31848
rect 24275 31808 24307 31816
tri 24307 31808 24315 31816 sw
tri 24393 31808 24401 31816 ne
rect 24401 31808 24455 31816
tri 24455 31808 24495 31848 sw
tri 24541 31808 24581 31848 ne
rect 24581 31830 24635 31848
tri 24635 31830 24653 31848 sw
tri 24721 31830 24739 31848 ne
rect 24739 31830 24815 31848
rect 24581 31822 24653 31830
tri 24653 31822 24661 31830 sw
tri 24739 31822 24747 31830 ne
rect 24747 31822 24815 31830
tri 24815 31822 24841 31848 sw
rect 24581 31808 24661 31822
tri 24661 31808 24675 31822 sw
tri 24747 31808 24761 31822 ne
rect 24761 31808 24841 31822
rect 24275 31754 24315 31808
tri 24315 31754 24369 31808 sw
tri 24401 31754 24455 31808 ne
rect 24455 31776 24495 31808
tri 24495 31776 24527 31808 sw
tri 24581 31776 24613 31808 ne
rect 24613 31776 24675 31808
rect 24455 31768 24527 31776
tri 24527 31768 24535 31776 sw
tri 24613 31768 24621 31776 ne
rect 24621 31768 24675 31776
tri 24675 31768 24715 31808 sw
tri 24761 31794 24775 31808 ne
rect 24455 31754 24535 31768
tri 24535 31754 24549 31768 sw
tri 24621 31754 24635 31768 ne
rect 24635 31754 24715 31768
tri 24275 31660 24369 31754 ne
tri 24369 31722 24401 31754 sw
tri 24455 31722 24487 31754 ne
rect 24487 31722 24549 31754
rect 24369 31714 24401 31722
tri 24401 31714 24409 31722 sw
tri 24487 31714 24495 31722 ne
rect 24495 31714 24549 31722
tri 24549 31714 24589 31754 sw
tri 24635 31740 24649 31754 ne
rect 24369 31660 24409 31714
tri 24409 31660 24463 31714 sw
tri 24495 31686 24523 31714 ne
tri 24369 31632 24397 31660 ne
rect 24397 29920 24463 31660
rect 24397 29864 24402 29920
rect 24458 29864 24463 29920
rect 24397 29840 24463 29864
rect 24397 29784 24402 29840
rect 24458 29784 24463 29840
rect 24397 29767 24463 29784
tri 5567 29493 5647 29573 sw
rect 5501 29488 5647 29493
rect 5501 29432 5506 29488
rect 5562 29432 5586 29488
rect 5642 29432 5647 29488
rect 5501 29427 5647 29432
rect 5295 29388 5441 29393
rect 5295 29332 5300 29388
rect 5356 29332 5380 29388
rect 5436 29332 5441 29388
rect 5295 29327 5441 29332
rect 21299 27345 21892 27790
rect 24523 21096 24589 31714
rect 24649 18589 24715 31754
rect 24775 20822 24841 31808
rect 24775 20766 24780 20822
rect 24836 20766 24841 20822
rect 24775 20742 24841 20766
rect 24775 20686 24780 20742
rect 24836 20686 24841 20742
rect 24775 20677 24841 20686
rect 24901 20105 24967 31862
rect 25027 21231 25093 31930
rect 25027 21175 25032 21231
rect 25088 21175 25093 21231
rect 25027 21151 25093 21175
rect 25027 21095 25032 21151
rect 25088 21095 25093 21151
rect 25027 21090 25093 21095
rect 25154 21137 25220 31984
rect 25154 21081 25159 21137
rect 25215 21081 25220 21137
rect 25154 21057 25220 21081
rect 25154 21001 25159 21057
rect 25215 21001 25220 21057
rect 25154 20996 25220 21001
rect 24901 20049 24906 20105
rect 24962 20049 24967 20105
rect 24901 20025 24967 20049
rect 24901 19969 24906 20025
rect 24962 19969 24967 20025
rect 24901 19960 24967 19969
rect 24649 18533 24654 18589
rect 24710 18533 24715 18589
rect 24649 18509 24715 18533
rect 2646 18462 2686 18491
rect 24649 18453 24654 18509
rect 24710 18453 24715 18509
rect 24649 18444 24715 18453
use sky130_fd_io__gpio_ovtv2_obpredrvr_new_i2c_fix_leak_fix  sky130_fd_io__gpio_ovtv2_obpredrvr_new_i2c_fix_leak_fix_0
timestamp 1683767628
transform 1 0 -49 0 1 28727
box 255 -19630 28132 5180
use sky130_fd_io__gpio_ovtv2_obpredrvr_old  sky130_fd_io__gpio_ovtv2_obpredrvr_old_0
timestamp 1683767628
transform 0 1 23158 -1 0 30683
box -255 631 13433 4925
<< labels >>
flabel metal3 s 2646 18462 2686 18491 0 FreeSans 200 0 0 0 NGHS_H
port 2 nsew
flabel metal3 s 21299 27345 21892 27790 3 FreeSans 520 270 0 0 VGND_IO
port 3 nsew
flabel metal3 s 21595 27567 21595 27567 3 FreeSans 520 270 0 0 VGND_IO
flabel metal1 s 11513 32365 11551 32404 3 FreeSans 520 90 0 0 OE_I_H_N
port 5 nsew
flabel metal1 s 26335 17905 26537 17947 7 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 25923 17881 26053 17923 7 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 25307 17775 25437 17817 7 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 24184 17775 24386 17817 7 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 24184 29706 24386 29748 3 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 25923 30641 26053 30683 3 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 26335 30641 26537 30683 3 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 26861 17775 27063 17817 7 FreeSans 300 270 0 0 VCC_IO
port 6 nsew
flabel metal1 s 27575 17775 27721 17812 7 FreeSans 300 270 0 0 VCC_IO
port 6 nsew
flabel metal1 s 24710 17775 24912 17817 7 FreeSans 300 270 0 0 VCC_IO
port 6 nsew
flabel metal1 s 24432 30637 24634 30679 3 FreeSans 300 270 0 0 VCC_IO
port 6 nsew
flabel metal1 s 27575 30646 27721 30683 3 FreeSans 300 270 0 0 VCC_IO
port 6 nsew
flabel metal1 s 26861 30641 27063 30683 3 FreeSans 300 270 0 0 VCC_IO
port 6 nsew
flabel metal1 s 25465 20856 25511 20902 3 FreeSans 300 270 0 0 SLOW_H
port 7 nsew
flabel metal1 s 27321 30418 27352 30562 3 FreeSans 520 270 0 0 PUEN_H[1]
port 8 nsew
flabel metal1 s 26721 23039 26752 23133 3 FreeSans 520 270 0 0 PUEN_H[0]
port 9 nsew
flabel metal1 s 27091 24740 27137 24781 3 FreeSans 300 270 0 0 PU_H_N[3]
port 10 nsew
flabel metal1 s 27091 24877 27137 24917 7 FreeSans 300 270 0 0 PU_H_N[2]
port 11 nsew
flabel metal1 s 27247 20545 27293 20585 3 FreeSans 300 270 0 0 PU_H_N[1]
port 12 nsew
flabel metal1 s 27171 22975 27217 23015 3 FreeSans 300 270 0 0 PU_H_N[0]
port 13 nsew
flabel metal1 s 27289 21535 27335 21581 3 FreeSans 300 270 0 0 PD_H[1]
port 14 nsew
flabel metal1 s 18581 32317 19176 32472 3 FreeSans 520 90 0 0 VGND_IO
port 3 nsew
flabel metal1 s 18522 33471 19108 33673 3 FreeSans 520 90 0 0 VCC_IO
port 6 nsew
flabel metal1 s 27289 22777 27335 22823 3 FreeSans 300 270 0 0 PD_H[0]
port 15 nsew
flabel metal1 s 26650 22321 26674 22407 3 FreeSans 520 270 0 0 PDEN_H_N[0]
port 16 nsew
flabel metal2 s 4839 28595 4994 28884 3 FreeSans 520 180 0 0 VGND_IO
port 3 nsew
flabel metal2 s 4916 28739 4916 28739 3 FreeSans 520 180 0 0 VGND_IO
flabel metal2 s 11274 33500 11643 33685 3 FreeSans 520 90 0 0 VCC_IO
port 6 nsew
flabel metal2 s 2028 29282 2200 29364 3 FreeSans 520 0 0 0 PD_H[3]
port 18 nsew
flabel metal2 s 2114 29323 2114 29323 3 FreeSans 520 0 0 0 PD_H[3]
flabel metal2 s 2214 29431 2333 29489 3 FreeSans 520 0 0 0 PD_H[2]
port 19 nsew
flabel metal2 s 18919 27043 19027 27411 3 FreeSans 520 180 0 0 PAD
port 20 nsew
flabel metal2 s 22701 27039 22809 27407 3 FreeSans 520 0 0 0 PAD
port 20 nsew
flabel metal2 s 22755 27223 22755 27223 3 FreeSans 520 0 0 0 PAD
flabel metal2 s 25722 23272 25873 23315 3 FreeSans 520 270 0 0 PDEN_H_N[1]
port 21 nsew
flabel metal2 s 26781 20301 26833 20359 3 FreeSans 300 270 0 0 PD_H[3]
port 18 nsew
flabel metal2 s 25098 20781 25150 20828 3 FreeSans 300 270 0 0 PD_H[2]
port 19 nsew
flabel metal2 s 26621 17940 26673 17987 7 FreeSans 300 270 0 0 DRVLO_H_N
port 22 nsew
flabel metal2 s 26693 23756 26745 23808 3 FreeSans 300 270 0 0 DRVHI_H
port 23 nsew
flabel locali s 18234 32803 18269 32838 3 FreeSans 520 90 0 0 SLOW_H_N
port 24 nsew
flabel locali s 19211 32744 19267 32788 3 FreeSans 520 90 0 0 SLEW_CTL_H_N[0]
port 25 nsew
flabel locali s 18420 32797 18456 32833 3 FreeSans 520 90 0 0 SLEW_CTL_H[1]
port 26 nsew
flabel locali s 16965 32758 16996 32798 3 FreeSans 520 90 0 0 PDEN_H_N[1]
port 21 nsew
flabel locali s 11923 32808 11954 32846 3 FreeSans 520 90 0 0 PD_DIS_H
port 27 nsew
flabel locali s 18056 32815 18086 32844 3 FreeSans 520 90 0 0 I2C_MODE_H_N
port 28 nsew
flabel locali s 16799 32751 16831 32795 3 FreeSans 520 90 0 0 DRVLO_H_N
port 22 nsew
<< properties >>
string GDS_END 38188490
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 38172632
<< end >>
