magic
tech sky130B
magscale 1 2
timestamp 1683767628
use sky130_fd_pr__dfl1sd2__example_5595914180884  sky130_fd_pr__dfl1sd2__example_5595914180884_0
timestamp 1683767628
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180884  sky130_fd_pr__dfl1sd2__example_5595914180884_1
timestamp 1683767628
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180884  sky130_fd_pr__dfl1sd2__example_5595914180884_2
timestamp 1683767628
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180884  sky130_fd_pr__dfl1sd2__example_5595914180884_3
timestamp 1683767628
transform 1 0 568 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180884  sky130_fd_pr__dfl1sd2__example_5595914180884_4
timestamp 1683767628
transform 1 0 724 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180819  sky130_fd_pr__dfl1sd__example_5595914180819_0
timestamp 1683767628
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180819  sky130_fd_pr__dfl1sd__example_5595914180819_1
timestamp 1683767628
transform 1 0 880 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 40073688
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 40070196
<< end >>
