magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -1396 -5168 1396 5168
<< pwell >>
rect -1962 5320 1962 5766
rect -1962 -5320 -1516 5320
rect 1516 -5320 1962 5320
rect -1962 -5766 1962 -5320
<< mvpsubdiff >>
rect -1936 5730 1936 5740
rect -1936 5356 -1411 5730
rect 1411 5356 1936 5730
rect -1936 5346 1936 5356
rect -1936 5219 -1542 5346
rect -1936 -5219 -1926 5219
rect -1552 -5219 -1542 5219
rect 1542 5219 1936 5346
rect -1936 -5346 -1542 -5219
rect 1542 -5219 1552 5219
rect 1926 -5219 1936 5219
rect 1542 -5346 1936 -5219
rect -1936 -5356 1936 -5346
rect -1936 -5730 -1411 -5356
rect 1411 -5730 1936 -5356
rect -1936 -5740 1936 -5730
<< mvnsubdiff >>
rect -1330 5068 -1183 5102
rect -1149 5068 -1115 5102
rect -1081 5068 -1047 5102
rect -1013 5068 -979 5102
rect -945 5068 -651 5102
rect -617 5068 -583 5102
rect -549 5068 -515 5102
rect -481 5068 -447 5102
rect -413 5068 -119 5102
rect -85 5068 -51 5102
rect -17 5068 17 5102
rect 51 5068 85 5102
rect 119 5068 413 5102
rect 447 5068 481 5102
rect 515 5068 549 5102
rect 583 5068 617 5102
rect 651 5068 945 5102
rect 979 5068 1013 5102
rect 1047 5068 1081 5102
rect 1115 5068 1149 5102
rect 1183 5068 1330 5102
rect -1330 5015 -1232 5068
rect -1330 4981 -1266 5015
rect -896 5015 -700 5068
rect -1330 4947 -1232 4981
rect -1330 4913 -1266 4947
rect -1330 4879 -1232 4913
rect -1330 4845 -1266 4879
rect -1330 4811 -1232 4845
rect -1330 4777 -1266 4811
rect -1330 4743 -1232 4777
rect -1330 4709 -1266 4743
rect -1330 4675 -1232 4709
rect -1330 4641 -1266 4675
rect -1330 4607 -1232 4641
rect -1330 4573 -1266 4607
rect -1330 4539 -1232 4573
rect -1330 4505 -1266 4539
rect -1330 4471 -1232 4505
rect -1330 4437 -1266 4471
rect -1330 4403 -1232 4437
rect -1330 4369 -1266 4403
rect -1330 4335 -1232 4369
rect -1330 4301 -1266 4335
rect -1330 4267 -1232 4301
rect -1330 4233 -1266 4267
rect -1330 4199 -1232 4233
rect -1330 4165 -1266 4199
rect -1330 4131 -1232 4165
rect -1330 4097 -1266 4131
rect -1330 4063 -1232 4097
rect -1330 4029 -1266 4063
rect -1330 3995 -1232 4029
rect -1330 3961 -1266 3995
rect -1330 3927 -1232 3961
rect -1330 3893 -1266 3927
rect -1330 3859 -1232 3893
rect -1330 3825 -1266 3859
rect -1330 3791 -1232 3825
rect -1330 3757 -1266 3791
rect -1330 3723 -1232 3757
rect -1330 3689 -1266 3723
rect -1330 3655 -1232 3689
rect -1330 3621 -1266 3655
rect -1330 3587 -1232 3621
rect -1330 3553 -1266 3587
rect -1330 3519 -1232 3553
rect -1330 3485 -1266 3519
rect -1330 3451 -1232 3485
rect -1330 3417 -1266 3451
rect -1330 3383 -1232 3417
rect -1330 3349 -1266 3383
rect -1330 3315 -1232 3349
rect -1330 3281 -1266 3315
rect -1330 3247 -1232 3281
rect -1330 3213 -1266 3247
rect -1330 3179 -1232 3213
rect -1330 3145 -1266 3179
rect -1330 3111 -1232 3145
rect -1330 3077 -1266 3111
rect -1330 3043 -1232 3077
rect -1330 3009 -1266 3043
rect -1330 2975 -1232 3009
rect -1330 2941 -1266 2975
rect -1330 2907 -1232 2941
rect -1330 2873 -1266 2907
rect -1330 2839 -1232 2873
rect -1330 2805 -1266 2839
rect -1330 2771 -1232 2805
rect -1330 2737 -1266 2771
rect -1330 2703 -1232 2737
rect -1330 2669 -1266 2703
rect -1330 2635 -1232 2669
rect -1330 2601 -1266 2635
rect -1330 2567 -1232 2601
rect -1330 2533 -1266 2567
rect -1330 2499 -1232 2533
rect -1330 2465 -1266 2499
rect -1330 2431 -1232 2465
rect -1330 2397 -1266 2431
rect -1330 2363 -1232 2397
rect -1330 2329 -1266 2363
rect -1330 2295 -1232 2329
rect -1330 2261 -1266 2295
rect -1330 2227 -1232 2261
rect -1330 2193 -1266 2227
rect -1330 2159 -1232 2193
rect -1330 2125 -1266 2159
rect -1330 2091 -1232 2125
rect -1330 2057 -1266 2091
rect -1330 2023 -1232 2057
rect -1330 1989 -1266 2023
rect -1330 1955 -1232 1989
rect -1330 1921 -1266 1955
rect -1330 1887 -1232 1921
rect -1330 1853 -1266 1887
rect -1330 1819 -1232 1853
rect -1330 1785 -1266 1819
rect -1330 1751 -1232 1785
rect -1330 1717 -1266 1751
rect -1330 1683 -1232 1717
rect -1330 1649 -1266 1683
rect -1330 1615 -1232 1649
rect -1330 1581 -1266 1615
rect -1330 1547 -1232 1581
rect -1330 1513 -1266 1547
rect -1330 1479 -1232 1513
rect -1330 1445 -1266 1479
rect -1330 1411 -1232 1445
rect -1330 1377 -1266 1411
rect -1330 1343 -1232 1377
rect -1330 1309 -1266 1343
rect -1330 1275 -1232 1309
rect -1330 1241 -1266 1275
rect -1330 1207 -1232 1241
rect -1330 1173 -1266 1207
rect -1330 1139 -1232 1173
rect -1330 1105 -1266 1139
rect -1330 1071 -1232 1105
rect -1330 1037 -1266 1071
rect -1330 1003 -1232 1037
rect -1330 969 -1266 1003
rect -1330 935 -1232 969
rect -1330 901 -1266 935
rect -1330 867 -1232 901
rect -1330 833 -1266 867
rect -1330 799 -1232 833
rect -1330 765 -1266 799
rect -1330 731 -1232 765
rect -1330 697 -1266 731
rect -1330 663 -1232 697
rect -1330 629 -1266 663
rect -1330 595 -1232 629
rect -1330 561 -1266 595
rect -1330 527 -1232 561
rect -1330 493 -1266 527
rect -1330 459 -1232 493
rect -1330 425 -1266 459
rect -1330 391 -1232 425
rect -1330 357 -1266 391
rect -1330 323 -1232 357
rect -1330 289 -1266 323
rect -1330 255 -1232 289
rect -1330 221 -1266 255
rect -1330 187 -1232 221
rect -1330 153 -1266 187
rect -1330 119 -1232 153
rect -1330 85 -1266 119
rect -1330 51 -1232 85
rect -1330 17 -1266 51
rect -1330 -17 -1232 17
rect -1330 -51 -1266 -17
rect -1330 -85 -1232 -51
rect -1330 -119 -1266 -85
rect -1330 -153 -1232 -119
rect -1330 -187 -1266 -153
rect -1330 -221 -1232 -187
rect -1330 -255 -1266 -221
rect -1330 -289 -1232 -255
rect -1330 -323 -1266 -289
rect -1330 -357 -1232 -323
rect -1330 -391 -1266 -357
rect -1330 -425 -1232 -391
rect -1330 -459 -1266 -425
rect -1330 -493 -1232 -459
rect -1330 -527 -1266 -493
rect -1330 -561 -1232 -527
rect -1330 -595 -1266 -561
rect -1330 -629 -1232 -595
rect -1330 -663 -1266 -629
rect -1330 -697 -1232 -663
rect -1330 -731 -1266 -697
rect -1330 -765 -1232 -731
rect -1330 -799 -1266 -765
rect -1330 -833 -1232 -799
rect -1330 -867 -1266 -833
rect -1330 -901 -1232 -867
rect -1330 -935 -1266 -901
rect -1330 -969 -1232 -935
rect -1330 -1003 -1266 -969
rect -1330 -1037 -1232 -1003
rect -1330 -1071 -1266 -1037
rect -1330 -1105 -1232 -1071
rect -1330 -1139 -1266 -1105
rect -1330 -1173 -1232 -1139
rect -1330 -1207 -1266 -1173
rect -1330 -1241 -1232 -1207
rect -1330 -1275 -1266 -1241
rect -1330 -1309 -1232 -1275
rect -1330 -1343 -1266 -1309
rect -1330 -1377 -1232 -1343
rect -1330 -1411 -1266 -1377
rect -1330 -1445 -1232 -1411
rect -1330 -1479 -1266 -1445
rect -1330 -1513 -1232 -1479
rect -1330 -1547 -1266 -1513
rect -1330 -1581 -1232 -1547
rect -1330 -1615 -1266 -1581
rect -1330 -1649 -1232 -1615
rect -1330 -1683 -1266 -1649
rect -1330 -1717 -1232 -1683
rect -1330 -1751 -1266 -1717
rect -1330 -1785 -1232 -1751
rect -1330 -1819 -1266 -1785
rect -1330 -1853 -1232 -1819
rect -1330 -1887 -1266 -1853
rect -1330 -1921 -1232 -1887
rect -1330 -1955 -1266 -1921
rect -1330 -1989 -1232 -1955
rect -1330 -2023 -1266 -1989
rect -1330 -2057 -1232 -2023
rect -1330 -2091 -1266 -2057
rect -1330 -2125 -1232 -2091
rect -1330 -2159 -1266 -2125
rect -1330 -2193 -1232 -2159
rect -1330 -2227 -1266 -2193
rect -1330 -2261 -1232 -2227
rect -1330 -2295 -1266 -2261
rect -1330 -2329 -1232 -2295
rect -1330 -2363 -1266 -2329
rect -1330 -2397 -1232 -2363
rect -1330 -2431 -1266 -2397
rect -1330 -2465 -1232 -2431
rect -1330 -2499 -1266 -2465
rect -1330 -2533 -1232 -2499
rect -1330 -2567 -1266 -2533
rect -1330 -2601 -1232 -2567
rect -1330 -2635 -1266 -2601
rect -1330 -2669 -1232 -2635
rect -1330 -2703 -1266 -2669
rect -1330 -2737 -1232 -2703
rect -1330 -2771 -1266 -2737
rect -1330 -2805 -1232 -2771
rect -1330 -2839 -1266 -2805
rect -1330 -2873 -1232 -2839
rect -1330 -2907 -1266 -2873
rect -1330 -2941 -1232 -2907
rect -1330 -2975 -1266 -2941
rect -1330 -3009 -1232 -2975
rect -1330 -3043 -1266 -3009
rect -1330 -3077 -1232 -3043
rect -1330 -3111 -1266 -3077
rect -1330 -3145 -1232 -3111
rect -1330 -3179 -1266 -3145
rect -1330 -3213 -1232 -3179
rect -1330 -3247 -1266 -3213
rect -1330 -3281 -1232 -3247
rect -1330 -3315 -1266 -3281
rect -1330 -3349 -1232 -3315
rect -1330 -3383 -1266 -3349
rect -1330 -3417 -1232 -3383
rect -1330 -3451 -1266 -3417
rect -1330 -3485 -1232 -3451
rect -1330 -3519 -1266 -3485
rect -1330 -3553 -1232 -3519
rect -1330 -3587 -1266 -3553
rect -1330 -3621 -1232 -3587
rect -1330 -3655 -1266 -3621
rect -1330 -3689 -1232 -3655
rect -1330 -3723 -1266 -3689
rect -1330 -3757 -1232 -3723
rect -1330 -3791 -1266 -3757
rect -1330 -3825 -1232 -3791
rect -1330 -3859 -1266 -3825
rect -1330 -3893 -1232 -3859
rect -1330 -3927 -1266 -3893
rect -1330 -3961 -1232 -3927
rect -1330 -3995 -1266 -3961
rect -1330 -4029 -1232 -3995
rect -1330 -4063 -1266 -4029
rect -1330 -4097 -1232 -4063
rect -1330 -4131 -1266 -4097
rect -1330 -4165 -1232 -4131
rect -1330 -4199 -1266 -4165
rect -1330 -4233 -1232 -4199
rect -1330 -4267 -1266 -4233
rect -1330 -4301 -1232 -4267
rect -1330 -4335 -1266 -4301
rect -1330 -4369 -1232 -4335
rect -1330 -4403 -1266 -4369
rect -1330 -4437 -1232 -4403
rect -1330 -4471 -1266 -4437
rect -1330 -4505 -1232 -4471
rect -1330 -4539 -1266 -4505
rect -1330 -4573 -1232 -4539
rect -1330 -4607 -1266 -4573
rect -1330 -4641 -1232 -4607
rect -1330 -4675 -1266 -4641
rect -1330 -4709 -1232 -4675
rect -1330 -4743 -1266 -4709
rect -1330 -4777 -1232 -4743
rect -1330 -4811 -1266 -4777
rect -1330 -4845 -1232 -4811
rect -1330 -4879 -1266 -4845
rect -1330 -4913 -1232 -4879
rect -1330 -4947 -1266 -4913
rect -1330 -4981 -1232 -4947
rect -1330 -5015 -1266 -4981
rect -862 4981 -815 5015
rect -781 4981 -734 5015
rect -364 5015 -168 5068
rect -896 4947 -700 4981
rect -862 4913 -815 4947
rect -781 4913 -734 4947
rect -896 4879 -700 4913
rect -862 4845 -815 4879
rect -781 4845 -734 4879
rect -896 4811 -700 4845
rect -862 4777 -815 4811
rect -781 4777 -734 4811
rect -896 4743 -700 4777
rect -862 4709 -815 4743
rect -781 4709 -734 4743
rect -896 4675 -700 4709
rect -862 4641 -815 4675
rect -781 4641 -734 4675
rect -896 4607 -700 4641
rect -862 4573 -815 4607
rect -781 4573 -734 4607
rect -896 4539 -700 4573
rect -862 4505 -815 4539
rect -781 4505 -734 4539
rect -896 4471 -700 4505
rect -862 4437 -815 4471
rect -781 4437 -734 4471
rect -896 4403 -700 4437
rect -862 4369 -815 4403
rect -781 4369 -734 4403
rect -896 4335 -700 4369
rect -862 4301 -815 4335
rect -781 4301 -734 4335
rect -896 4267 -700 4301
rect -862 4233 -815 4267
rect -781 4233 -734 4267
rect -896 4199 -700 4233
rect -862 4165 -815 4199
rect -781 4165 -734 4199
rect -896 4131 -700 4165
rect -862 4097 -815 4131
rect -781 4097 -734 4131
rect -896 4063 -700 4097
rect -862 4029 -815 4063
rect -781 4029 -734 4063
rect -896 3995 -700 4029
rect -862 3961 -815 3995
rect -781 3961 -734 3995
rect -896 3927 -700 3961
rect -862 3893 -815 3927
rect -781 3893 -734 3927
rect -896 3859 -700 3893
rect -862 3825 -815 3859
rect -781 3825 -734 3859
rect -896 3791 -700 3825
rect -862 3757 -815 3791
rect -781 3757 -734 3791
rect -896 3723 -700 3757
rect -862 3689 -815 3723
rect -781 3689 -734 3723
rect -896 3655 -700 3689
rect -862 3621 -815 3655
rect -781 3621 -734 3655
rect -896 3587 -700 3621
rect -862 3553 -815 3587
rect -781 3553 -734 3587
rect -896 3519 -700 3553
rect -862 3485 -815 3519
rect -781 3485 -734 3519
rect -896 3451 -700 3485
rect -862 3417 -815 3451
rect -781 3417 -734 3451
rect -896 3383 -700 3417
rect -862 3349 -815 3383
rect -781 3349 -734 3383
rect -896 3315 -700 3349
rect -862 3281 -815 3315
rect -781 3281 -734 3315
rect -896 3247 -700 3281
rect -862 3213 -815 3247
rect -781 3213 -734 3247
rect -896 3179 -700 3213
rect -862 3145 -815 3179
rect -781 3145 -734 3179
rect -896 3111 -700 3145
rect -862 3077 -815 3111
rect -781 3077 -734 3111
rect -896 3043 -700 3077
rect -862 3009 -815 3043
rect -781 3009 -734 3043
rect -896 2975 -700 3009
rect -862 2941 -815 2975
rect -781 2941 -734 2975
rect -896 2907 -700 2941
rect -862 2873 -815 2907
rect -781 2873 -734 2907
rect -896 2839 -700 2873
rect -862 2805 -815 2839
rect -781 2805 -734 2839
rect -896 2771 -700 2805
rect -862 2737 -815 2771
rect -781 2737 -734 2771
rect -896 2703 -700 2737
rect -862 2669 -815 2703
rect -781 2669 -734 2703
rect -896 2635 -700 2669
rect -862 2601 -815 2635
rect -781 2601 -734 2635
rect -896 2567 -700 2601
rect -862 2533 -815 2567
rect -781 2533 -734 2567
rect -896 2499 -700 2533
rect -862 2465 -815 2499
rect -781 2465 -734 2499
rect -896 2431 -700 2465
rect -862 2397 -815 2431
rect -781 2397 -734 2431
rect -896 2363 -700 2397
rect -862 2329 -815 2363
rect -781 2329 -734 2363
rect -896 2295 -700 2329
rect -862 2261 -815 2295
rect -781 2261 -734 2295
rect -896 2227 -700 2261
rect -862 2193 -815 2227
rect -781 2193 -734 2227
rect -896 2159 -700 2193
rect -862 2125 -815 2159
rect -781 2125 -734 2159
rect -896 2091 -700 2125
rect -862 2057 -815 2091
rect -781 2057 -734 2091
rect -896 2023 -700 2057
rect -862 1989 -815 2023
rect -781 1989 -734 2023
rect -896 1955 -700 1989
rect -862 1921 -815 1955
rect -781 1921 -734 1955
rect -896 1887 -700 1921
rect -862 1853 -815 1887
rect -781 1853 -734 1887
rect -896 1819 -700 1853
rect -862 1785 -815 1819
rect -781 1785 -734 1819
rect -896 1751 -700 1785
rect -862 1717 -815 1751
rect -781 1717 -734 1751
rect -896 1683 -700 1717
rect -862 1649 -815 1683
rect -781 1649 -734 1683
rect -896 1615 -700 1649
rect -862 1581 -815 1615
rect -781 1581 -734 1615
rect -896 1547 -700 1581
rect -862 1513 -815 1547
rect -781 1513 -734 1547
rect -896 1479 -700 1513
rect -862 1445 -815 1479
rect -781 1445 -734 1479
rect -896 1411 -700 1445
rect -862 1377 -815 1411
rect -781 1377 -734 1411
rect -896 1343 -700 1377
rect -862 1309 -815 1343
rect -781 1309 -734 1343
rect -896 1275 -700 1309
rect -862 1241 -815 1275
rect -781 1241 -734 1275
rect -896 1207 -700 1241
rect -862 1173 -815 1207
rect -781 1173 -734 1207
rect -896 1139 -700 1173
rect -862 1105 -815 1139
rect -781 1105 -734 1139
rect -896 1071 -700 1105
rect -862 1037 -815 1071
rect -781 1037 -734 1071
rect -896 1003 -700 1037
rect -862 969 -815 1003
rect -781 969 -734 1003
rect -896 935 -700 969
rect -862 901 -815 935
rect -781 901 -734 935
rect -896 867 -700 901
rect -862 833 -815 867
rect -781 833 -734 867
rect -896 799 -700 833
rect -862 765 -815 799
rect -781 765 -734 799
rect -896 731 -700 765
rect -862 697 -815 731
rect -781 697 -734 731
rect -896 663 -700 697
rect -862 629 -815 663
rect -781 629 -734 663
rect -896 595 -700 629
rect -862 561 -815 595
rect -781 561 -734 595
rect -896 527 -700 561
rect -862 493 -815 527
rect -781 493 -734 527
rect -896 459 -700 493
rect -862 425 -815 459
rect -781 425 -734 459
rect -896 391 -700 425
rect -862 357 -815 391
rect -781 357 -734 391
rect -896 323 -700 357
rect -862 289 -815 323
rect -781 289 -734 323
rect -896 255 -700 289
rect -862 221 -815 255
rect -781 221 -734 255
rect -896 187 -700 221
rect -862 153 -815 187
rect -781 153 -734 187
rect -896 119 -700 153
rect -862 85 -815 119
rect -781 85 -734 119
rect -896 51 -700 85
rect -862 17 -815 51
rect -781 17 -734 51
rect -896 -17 -700 17
rect -862 -51 -815 -17
rect -781 -51 -734 -17
rect -896 -85 -700 -51
rect -862 -119 -815 -85
rect -781 -119 -734 -85
rect -896 -153 -700 -119
rect -862 -187 -815 -153
rect -781 -187 -734 -153
rect -896 -221 -700 -187
rect -862 -255 -815 -221
rect -781 -255 -734 -221
rect -896 -289 -700 -255
rect -862 -323 -815 -289
rect -781 -323 -734 -289
rect -896 -357 -700 -323
rect -862 -391 -815 -357
rect -781 -391 -734 -357
rect -896 -425 -700 -391
rect -862 -459 -815 -425
rect -781 -459 -734 -425
rect -896 -493 -700 -459
rect -862 -527 -815 -493
rect -781 -527 -734 -493
rect -896 -561 -700 -527
rect -862 -595 -815 -561
rect -781 -595 -734 -561
rect -896 -629 -700 -595
rect -862 -663 -815 -629
rect -781 -663 -734 -629
rect -896 -697 -700 -663
rect -862 -731 -815 -697
rect -781 -731 -734 -697
rect -896 -765 -700 -731
rect -862 -799 -815 -765
rect -781 -799 -734 -765
rect -896 -833 -700 -799
rect -862 -867 -815 -833
rect -781 -867 -734 -833
rect -896 -901 -700 -867
rect -862 -935 -815 -901
rect -781 -935 -734 -901
rect -896 -969 -700 -935
rect -862 -1003 -815 -969
rect -781 -1003 -734 -969
rect -896 -1037 -700 -1003
rect -862 -1071 -815 -1037
rect -781 -1071 -734 -1037
rect -896 -1105 -700 -1071
rect -862 -1139 -815 -1105
rect -781 -1139 -734 -1105
rect -896 -1173 -700 -1139
rect -862 -1207 -815 -1173
rect -781 -1207 -734 -1173
rect -896 -1241 -700 -1207
rect -862 -1275 -815 -1241
rect -781 -1275 -734 -1241
rect -896 -1309 -700 -1275
rect -862 -1343 -815 -1309
rect -781 -1343 -734 -1309
rect -896 -1377 -700 -1343
rect -862 -1411 -815 -1377
rect -781 -1411 -734 -1377
rect -896 -1445 -700 -1411
rect -862 -1479 -815 -1445
rect -781 -1479 -734 -1445
rect -896 -1513 -700 -1479
rect -862 -1547 -815 -1513
rect -781 -1547 -734 -1513
rect -896 -1581 -700 -1547
rect -862 -1615 -815 -1581
rect -781 -1615 -734 -1581
rect -896 -1649 -700 -1615
rect -862 -1683 -815 -1649
rect -781 -1683 -734 -1649
rect -896 -1717 -700 -1683
rect -862 -1751 -815 -1717
rect -781 -1751 -734 -1717
rect -896 -1785 -700 -1751
rect -862 -1819 -815 -1785
rect -781 -1819 -734 -1785
rect -896 -1853 -700 -1819
rect -862 -1887 -815 -1853
rect -781 -1887 -734 -1853
rect -896 -1921 -700 -1887
rect -862 -1955 -815 -1921
rect -781 -1955 -734 -1921
rect -896 -1989 -700 -1955
rect -862 -2023 -815 -1989
rect -781 -2023 -734 -1989
rect -896 -2057 -700 -2023
rect -862 -2091 -815 -2057
rect -781 -2091 -734 -2057
rect -896 -2125 -700 -2091
rect -862 -2159 -815 -2125
rect -781 -2159 -734 -2125
rect -896 -2193 -700 -2159
rect -862 -2227 -815 -2193
rect -781 -2227 -734 -2193
rect -896 -2261 -700 -2227
rect -862 -2295 -815 -2261
rect -781 -2295 -734 -2261
rect -896 -2329 -700 -2295
rect -862 -2363 -815 -2329
rect -781 -2363 -734 -2329
rect -896 -2397 -700 -2363
rect -862 -2431 -815 -2397
rect -781 -2431 -734 -2397
rect -896 -2465 -700 -2431
rect -862 -2499 -815 -2465
rect -781 -2499 -734 -2465
rect -896 -2533 -700 -2499
rect -862 -2567 -815 -2533
rect -781 -2567 -734 -2533
rect -896 -2601 -700 -2567
rect -862 -2635 -815 -2601
rect -781 -2635 -734 -2601
rect -896 -2669 -700 -2635
rect -862 -2703 -815 -2669
rect -781 -2703 -734 -2669
rect -896 -2737 -700 -2703
rect -862 -2771 -815 -2737
rect -781 -2771 -734 -2737
rect -896 -2805 -700 -2771
rect -862 -2839 -815 -2805
rect -781 -2839 -734 -2805
rect -896 -2873 -700 -2839
rect -862 -2907 -815 -2873
rect -781 -2907 -734 -2873
rect -896 -2941 -700 -2907
rect -862 -2975 -815 -2941
rect -781 -2975 -734 -2941
rect -896 -3009 -700 -2975
rect -862 -3043 -815 -3009
rect -781 -3043 -734 -3009
rect -896 -3077 -700 -3043
rect -862 -3111 -815 -3077
rect -781 -3111 -734 -3077
rect -896 -3145 -700 -3111
rect -862 -3179 -815 -3145
rect -781 -3179 -734 -3145
rect -896 -3213 -700 -3179
rect -862 -3247 -815 -3213
rect -781 -3247 -734 -3213
rect -896 -3281 -700 -3247
rect -862 -3315 -815 -3281
rect -781 -3315 -734 -3281
rect -896 -3349 -700 -3315
rect -862 -3383 -815 -3349
rect -781 -3383 -734 -3349
rect -896 -3417 -700 -3383
rect -862 -3451 -815 -3417
rect -781 -3451 -734 -3417
rect -896 -3485 -700 -3451
rect -862 -3519 -815 -3485
rect -781 -3519 -734 -3485
rect -896 -3553 -700 -3519
rect -862 -3587 -815 -3553
rect -781 -3587 -734 -3553
rect -896 -3621 -700 -3587
rect -862 -3655 -815 -3621
rect -781 -3655 -734 -3621
rect -896 -3689 -700 -3655
rect -862 -3723 -815 -3689
rect -781 -3723 -734 -3689
rect -896 -3757 -700 -3723
rect -862 -3791 -815 -3757
rect -781 -3791 -734 -3757
rect -896 -3825 -700 -3791
rect -862 -3859 -815 -3825
rect -781 -3859 -734 -3825
rect -896 -3893 -700 -3859
rect -862 -3927 -815 -3893
rect -781 -3927 -734 -3893
rect -896 -3961 -700 -3927
rect -862 -3995 -815 -3961
rect -781 -3995 -734 -3961
rect -896 -4029 -700 -3995
rect -862 -4063 -815 -4029
rect -781 -4063 -734 -4029
rect -896 -4097 -700 -4063
rect -862 -4131 -815 -4097
rect -781 -4131 -734 -4097
rect -896 -4165 -700 -4131
rect -862 -4199 -815 -4165
rect -781 -4199 -734 -4165
rect -896 -4233 -700 -4199
rect -862 -4267 -815 -4233
rect -781 -4267 -734 -4233
rect -896 -4301 -700 -4267
rect -862 -4335 -815 -4301
rect -781 -4335 -734 -4301
rect -896 -4369 -700 -4335
rect -862 -4403 -815 -4369
rect -781 -4403 -734 -4369
rect -896 -4437 -700 -4403
rect -862 -4471 -815 -4437
rect -781 -4471 -734 -4437
rect -896 -4505 -700 -4471
rect -862 -4539 -815 -4505
rect -781 -4539 -734 -4505
rect -896 -4573 -700 -4539
rect -862 -4607 -815 -4573
rect -781 -4607 -734 -4573
rect -896 -4641 -700 -4607
rect -862 -4675 -815 -4641
rect -781 -4675 -734 -4641
rect -896 -4709 -700 -4675
rect -862 -4743 -815 -4709
rect -781 -4743 -734 -4709
rect -896 -4777 -700 -4743
rect -862 -4811 -815 -4777
rect -781 -4811 -734 -4777
rect -896 -4845 -700 -4811
rect -862 -4879 -815 -4845
rect -781 -4879 -734 -4845
rect -896 -4913 -700 -4879
rect -862 -4947 -815 -4913
rect -781 -4947 -734 -4913
rect -896 -4981 -700 -4947
rect -1330 -5068 -1232 -5015
rect -862 -5015 -815 -4981
rect -781 -5015 -734 -4981
rect -330 4981 -283 5015
rect -249 4981 -202 5015
rect 168 5015 364 5068
rect -364 4947 -168 4981
rect -330 4913 -283 4947
rect -249 4913 -202 4947
rect -364 4879 -168 4913
rect -330 4845 -283 4879
rect -249 4845 -202 4879
rect -364 4811 -168 4845
rect -330 4777 -283 4811
rect -249 4777 -202 4811
rect -364 4743 -168 4777
rect -330 4709 -283 4743
rect -249 4709 -202 4743
rect -364 4675 -168 4709
rect -330 4641 -283 4675
rect -249 4641 -202 4675
rect -364 4607 -168 4641
rect -330 4573 -283 4607
rect -249 4573 -202 4607
rect -364 4539 -168 4573
rect -330 4505 -283 4539
rect -249 4505 -202 4539
rect -364 4471 -168 4505
rect -330 4437 -283 4471
rect -249 4437 -202 4471
rect -364 4403 -168 4437
rect -330 4369 -283 4403
rect -249 4369 -202 4403
rect -364 4335 -168 4369
rect -330 4301 -283 4335
rect -249 4301 -202 4335
rect -364 4267 -168 4301
rect -330 4233 -283 4267
rect -249 4233 -202 4267
rect -364 4199 -168 4233
rect -330 4165 -283 4199
rect -249 4165 -202 4199
rect -364 4131 -168 4165
rect -330 4097 -283 4131
rect -249 4097 -202 4131
rect -364 4063 -168 4097
rect -330 4029 -283 4063
rect -249 4029 -202 4063
rect -364 3995 -168 4029
rect -330 3961 -283 3995
rect -249 3961 -202 3995
rect -364 3927 -168 3961
rect -330 3893 -283 3927
rect -249 3893 -202 3927
rect -364 3859 -168 3893
rect -330 3825 -283 3859
rect -249 3825 -202 3859
rect -364 3791 -168 3825
rect -330 3757 -283 3791
rect -249 3757 -202 3791
rect -364 3723 -168 3757
rect -330 3689 -283 3723
rect -249 3689 -202 3723
rect -364 3655 -168 3689
rect -330 3621 -283 3655
rect -249 3621 -202 3655
rect -364 3587 -168 3621
rect -330 3553 -283 3587
rect -249 3553 -202 3587
rect -364 3519 -168 3553
rect -330 3485 -283 3519
rect -249 3485 -202 3519
rect -364 3451 -168 3485
rect -330 3417 -283 3451
rect -249 3417 -202 3451
rect -364 3383 -168 3417
rect -330 3349 -283 3383
rect -249 3349 -202 3383
rect -364 3315 -168 3349
rect -330 3281 -283 3315
rect -249 3281 -202 3315
rect -364 3247 -168 3281
rect -330 3213 -283 3247
rect -249 3213 -202 3247
rect -364 3179 -168 3213
rect -330 3145 -283 3179
rect -249 3145 -202 3179
rect -364 3111 -168 3145
rect -330 3077 -283 3111
rect -249 3077 -202 3111
rect -364 3043 -168 3077
rect -330 3009 -283 3043
rect -249 3009 -202 3043
rect -364 2975 -168 3009
rect -330 2941 -283 2975
rect -249 2941 -202 2975
rect -364 2907 -168 2941
rect -330 2873 -283 2907
rect -249 2873 -202 2907
rect -364 2839 -168 2873
rect -330 2805 -283 2839
rect -249 2805 -202 2839
rect -364 2771 -168 2805
rect -330 2737 -283 2771
rect -249 2737 -202 2771
rect -364 2703 -168 2737
rect -330 2669 -283 2703
rect -249 2669 -202 2703
rect -364 2635 -168 2669
rect -330 2601 -283 2635
rect -249 2601 -202 2635
rect -364 2567 -168 2601
rect -330 2533 -283 2567
rect -249 2533 -202 2567
rect -364 2499 -168 2533
rect -330 2465 -283 2499
rect -249 2465 -202 2499
rect -364 2431 -168 2465
rect -330 2397 -283 2431
rect -249 2397 -202 2431
rect -364 2363 -168 2397
rect -330 2329 -283 2363
rect -249 2329 -202 2363
rect -364 2295 -168 2329
rect -330 2261 -283 2295
rect -249 2261 -202 2295
rect -364 2227 -168 2261
rect -330 2193 -283 2227
rect -249 2193 -202 2227
rect -364 2159 -168 2193
rect -330 2125 -283 2159
rect -249 2125 -202 2159
rect -364 2091 -168 2125
rect -330 2057 -283 2091
rect -249 2057 -202 2091
rect -364 2023 -168 2057
rect -330 1989 -283 2023
rect -249 1989 -202 2023
rect -364 1955 -168 1989
rect -330 1921 -283 1955
rect -249 1921 -202 1955
rect -364 1887 -168 1921
rect -330 1853 -283 1887
rect -249 1853 -202 1887
rect -364 1819 -168 1853
rect -330 1785 -283 1819
rect -249 1785 -202 1819
rect -364 1751 -168 1785
rect -330 1717 -283 1751
rect -249 1717 -202 1751
rect -364 1683 -168 1717
rect -330 1649 -283 1683
rect -249 1649 -202 1683
rect -364 1615 -168 1649
rect -330 1581 -283 1615
rect -249 1581 -202 1615
rect -364 1547 -168 1581
rect -330 1513 -283 1547
rect -249 1513 -202 1547
rect -364 1479 -168 1513
rect -330 1445 -283 1479
rect -249 1445 -202 1479
rect -364 1411 -168 1445
rect -330 1377 -283 1411
rect -249 1377 -202 1411
rect -364 1343 -168 1377
rect -330 1309 -283 1343
rect -249 1309 -202 1343
rect -364 1275 -168 1309
rect -330 1241 -283 1275
rect -249 1241 -202 1275
rect -364 1207 -168 1241
rect -330 1173 -283 1207
rect -249 1173 -202 1207
rect -364 1139 -168 1173
rect -330 1105 -283 1139
rect -249 1105 -202 1139
rect -364 1071 -168 1105
rect -330 1037 -283 1071
rect -249 1037 -202 1071
rect -364 1003 -168 1037
rect -330 969 -283 1003
rect -249 969 -202 1003
rect -364 935 -168 969
rect -330 901 -283 935
rect -249 901 -202 935
rect -364 867 -168 901
rect -330 833 -283 867
rect -249 833 -202 867
rect -364 799 -168 833
rect -330 765 -283 799
rect -249 765 -202 799
rect -364 731 -168 765
rect -330 697 -283 731
rect -249 697 -202 731
rect -364 663 -168 697
rect -330 629 -283 663
rect -249 629 -202 663
rect -364 595 -168 629
rect -330 561 -283 595
rect -249 561 -202 595
rect -364 527 -168 561
rect -330 493 -283 527
rect -249 493 -202 527
rect -364 459 -168 493
rect -330 425 -283 459
rect -249 425 -202 459
rect -364 391 -168 425
rect -330 357 -283 391
rect -249 357 -202 391
rect -364 323 -168 357
rect -330 289 -283 323
rect -249 289 -202 323
rect -364 255 -168 289
rect -330 221 -283 255
rect -249 221 -202 255
rect -364 187 -168 221
rect -330 153 -283 187
rect -249 153 -202 187
rect -364 119 -168 153
rect -330 85 -283 119
rect -249 85 -202 119
rect -364 51 -168 85
rect -330 17 -283 51
rect -249 17 -202 51
rect -364 -17 -168 17
rect -330 -51 -283 -17
rect -249 -51 -202 -17
rect -364 -85 -168 -51
rect -330 -119 -283 -85
rect -249 -119 -202 -85
rect -364 -153 -168 -119
rect -330 -187 -283 -153
rect -249 -187 -202 -153
rect -364 -221 -168 -187
rect -330 -255 -283 -221
rect -249 -255 -202 -221
rect -364 -289 -168 -255
rect -330 -323 -283 -289
rect -249 -323 -202 -289
rect -364 -357 -168 -323
rect -330 -391 -283 -357
rect -249 -391 -202 -357
rect -364 -425 -168 -391
rect -330 -459 -283 -425
rect -249 -459 -202 -425
rect -364 -493 -168 -459
rect -330 -527 -283 -493
rect -249 -527 -202 -493
rect -364 -561 -168 -527
rect -330 -595 -283 -561
rect -249 -595 -202 -561
rect -364 -629 -168 -595
rect -330 -663 -283 -629
rect -249 -663 -202 -629
rect -364 -697 -168 -663
rect -330 -731 -283 -697
rect -249 -731 -202 -697
rect -364 -765 -168 -731
rect -330 -799 -283 -765
rect -249 -799 -202 -765
rect -364 -833 -168 -799
rect -330 -867 -283 -833
rect -249 -867 -202 -833
rect -364 -901 -168 -867
rect -330 -935 -283 -901
rect -249 -935 -202 -901
rect -364 -969 -168 -935
rect -330 -1003 -283 -969
rect -249 -1003 -202 -969
rect -364 -1037 -168 -1003
rect -330 -1071 -283 -1037
rect -249 -1071 -202 -1037
rect -364 -1105 -168 -1071
rect -330 -1139 -283 -1105
rect -249 -1139 -202 -1105
rect -364 -1173 -168 -1139
rect -330 -1207 -283 -1173
rect -249 -1207 -202 -1173
rect -364 -1241 -168 -1207
rect -330 -1275 -283 -1241
rect -249 -1275 -202 -1241
rect -364 -1309 -168 -1275
rect -330 -1343 -283 -1309
rect -249 -1343 -202 -1309
rect -364 -1377 -168 -1343
rect -330 -1411 -283 -1377
rect -249 -1411 -202 -1377
rect -364 -1445 -168 -1411
rect -330 -1479 -283 -1445
rect -249 -1479 -202 -1445
rect -364 -1513 -168 -1479
rect -330 -1547 -283 -1513
rect -249 -1547 -202 -1513
rect -364 -1581 -168 -1547
rect -330 -1615 -283 -1581
rect -249 -1615 -202 -1581
rect -364 -1649 -168 -1615
rect -330 -1683 -283 -1649
rect -249 -1683 -202 -1649
rect -364 -1717 -168 -1683
rect -330 -1751 -283 -1717
rect -249 -1751 -202 -1717
rect -364 -1785 -168 -1751
rect -330 -1819 -283 -1785
rect -249 -1819 -202 -1785
rect -364 -1853 -168 -1819
rect -330 -1887 -283 -1853
rect -249 -1887 -202 -1853
rect -364 -1921 -168 -1887
rect -330 -1955 -283 -1921
rect -249 -1955 -202 -1921
rect -364 -1989 -168 -1955
rect -330 -2023 -283 -1989
rect -249 -2023 -202 -1989
rect -364 -2057 -168 -2023
rect -330 -2091 -283 -2057
rect -249 -2091 -202 -2057
rect -364 -2125 -168 -2091
rect -330 -2159 -283 -2125
rect -249 -2159 -202 -2125
rect -364 -2193 -168 -2159
rect -330 -2227 -283 -2193
rect -249 -2227 -202 -2193
rect -364 -2261 -168 -2227
rect -330 -2295 -283 -2261
rect -249 -2295 -202 -2261
rect -364 -2329 -168 -2295
rect -330 -2363 -283 -2329
rect -249 -2363 -202 -2329
rect -364 -2397 -168 -2363
rect -330 -2431 -283 -2397
rect -249 -2431 -202 -2397
rect -364 -2465 -168 -2431
rect -330 -2499 -283 -2465
rect -249 -2499 -202 -2465
rect -364 -2533 -168 -2499
rect -330 -2567 -283 -2533
rect -249 -2567 -202 -2533
rect -364 -2601 -168 -2567
rect -330 -2635 -283 -2601
rect -249 -2635 -202 -2601
rect -364 -2669 -168 -2635
rect -330 -2703 -283 -2669
rect -249 -2703 -202 -2669
rect -364 -2737 -168 -2703
rect -330 -2771 -283 -2737
rect -249 -2771 -202 -2737
rect -364 -2805 -168 -2771
rect -330 -2839 -283 -2805
rect -249 -2839 -202 -2805
rect -364 -2873 -168 -2839
rect -330 -2907 -283 -2873
rect -249 -2907 -202 -2873
rect -364 -2941 -168 -2907
rect -330 -2975 -283 -2941
rect -249 -2975 -202 -2941
rect -364 -3009 -168 -2975
rect -330 -3043 -283 -3009
rect -249 -3043 -202 -3009
rect -364 -3077 -168 -3043
rect -330 -3111 -283 -3077
rect -249 -3111 -202 -3077
rect -364 -3145 -168 -3111
rect -330 -3179 -283 -3145
rect -249 -3179 -202 -3145
rect -364 -3213 -168 -3179
rect -330 -3247 -283 -3213
rect -249 -3247 -202 -3213
rect -364 -3281 -168 -3247
rect -330 -3315 -283 -3281
rect -249 -3315 -202 -3281
rect -364 -3349 -168 -3315
rect -330 -3383 -283 -3349
rect -249 -3383 -202 -3349
rect -364 -3417 -168 -3383
rect -330 -3451 -283 -3417
rect -249 -3451 -202 -3417
rect -364 -3485 -168 -3451
rect -330 -3519 -283 -3485
rect -249 -3519 -202 -3485
rect -364 -3553 -168 -3519
rect -330 -3587 -283 -3553
rect -249 -3587 -202 -3553
rect -364 -3621 -168 -3587
rect -330 -3655 -283 -3621
rect -249 -3655 -202 -3621
rect -364 -3689 -168 -3655
rect -330 -3723 -283 -3689
rect -249 -3723 -202 -3689
rect -364 -3757 -168 -3723
rect -330 -3791 -283 -3757
rect -249 -3791 -202 -3757
rect -364 -3825 -168 -3791
rect -330 -3859 -283 -3825
rect -249 -3859 -202 -3825
rect -364 -3893 -168 -3859
rect -330 -3927 -283 -3893
rect -249 -3927 -202 -3893
rect -364 -3961 -168 -3927
rect -330 -3995 -283 -3961
rect -249 -3995 -202 -3961
rect -364 -4029 -168 -3995
rect -330 -4063 -283 -4029
rect -249 -4063 -202 -4029
rect -364 -4097 -168 -4063
rect -330 -4131 -283 -4097
rect -249 -4131 -202 -4097
rect -364 -4165 -168 -4131
rect -330 -4199 -283 -4165
rect -249 -4199 -202 -4165
rect -364 -4233 -168 -4199
rect -330 -4267 -283 -4233
rect -249 -4267 -202 -4233
rect -364 -4301 -168 -4267
rect -330 -4335 -283 -4301
rect -249 -4335 -202 -4301
rect -364 -4369 -168 -4335
rect -330 -4403 -283 -4369
rect -249 -4403 -202 -4369
rect -364 -4437 -168 -4403
rect -330 -4471 -283 -4437
rect -249 -4471 -202 -4437
rect -364 -4505 -168 -4471
rect -330 -4539 -283 -4505
rect -249 -4539 -202 -4505
rect -364 -4573 -168 -4539
rect -330 -4607 -283 -4573
rect -249 -4607 -202 -4573
rect -364 -4641 -168 -4607
rect -330 -4675 -283 -4641
rect -249 -4675 -202 -4641
rect -364 -4709 -168 -4675
rect -330 -4743 -283 -4709
rect -249 -4743 -202 -4709
rect -364 -4777 -168 -4743
rect -330 -4811 -283 -4777
rect -249 -4811 -202 -4777
rect -364 -4845 -168 -4811
rect -330 -4879 -283 -4845
rect -249 -4879 -202 -4845
rect -364 -4913 -168 -4879
rect -330 -4947 -283 -4913
rect -249 -4947 -202 -4913
rect -364 -4981 -168 -4947
rect -896 -5068 -700 -5015
rect -330 -5015 -283 -4981
rect -249 -5015 -202 -4981
rect 202 4981 249 5015
rect 283 4981 330 5015
rect 700 5015 896 5068
rect 168 4947 364 4981
rect 202 4913 249 4947
rect 283 4913 330 4947
rect 168 4879 364 4913
rect 202 4845 249 4879
rect 283 4845 330 4879
rect 168 4811 364 4845
rect 202 4777 249 4811
rect 283 4777 330 4811
rect 168 4743 364 4777
rect 202 4709 249 4743
rect 283 4709 330 4743
rect 168 4675 364 4709
rect 202 4641 249 4675
rect 283 4641 330 4675
rect 168 4607 364 4641
rect 202 4573 249 4607
rect 283 4573 330 4607
rect 168 4539 364 4573
rect 202 4505 249 4539
rect 283 4505 330 4539
rect 168 4471 364 4505
rect 202 4437 249 4471
rect 283 4437 330 4471
rect 168 4403 364 4437
rect 202 4369 249 4403
rect 283 4369 330 4403
rect 168 4335 364 4369
rect 202 4301 249 4335
rect 283 4301 330 4335
rect 168 4267 364 4301
rect 202 4233 249 4267
rect 283 4233 330 4267
rect 168 4199 364 4233
rect 202 4165 249 4199
rect 283 4165 330 4199
rect 168 4131 364 4165
rect 202 4097 249 4131
rect 283 4097 330 4131
rect 168 4063 364 4097
rect 202 4029 249 4063
rect 283 4029 330 4063
rect 168 3995 364 4029
rect 202 3961 249 3995
rect 283 3961 330 3995
rect 168 3927 364 3961
rect 202 3893 249 3927
rect 283 3893 330 3927
rect 168 3859 364 3893
rect 202 3825 249 3859
rect 283 3825 330 3859
rect 168 3791 364 3825
rect 202 3757 249 3791
rect 283 3757 330 3791
rect 168 3723 364 3757
rect 202 3689 249 3723
rect 283 3689 330 3723
rect 168 3655 364 3689
rect 202 3621 249 3655
rect 283 3621 330 3655
rect 168 3587 364 3621
rect 202 3553 249 3587
rect 283 3553 330 3587
rect 168 3519 364 3553
rect 202 3485 249 3519
rect 283 3485 330 3519
rect 168 3451 364 3485
rect 202 3417 249 3451
rect 283 3417 330 3451
rect 168 3383 364 3417
rect 202 3349 249 3383
rect 283 3349 330 3383
rect 168 3315 364 3349
rect 202 3281 249 3315
rect 283 3281 330 3315
rect 168 3247 364 3281
rect 202 3213 249 3247
rect 283 3213 330 3247
rect 168 3179 364 3213
rect 202 3145 249 3179
rect 283 3145 330 3179
rect 168 3111 364 3145
rect 202 3077 249 3111
rect 283 3077 330 3111
rect 168 3043 364 3077
rect 202 3009 249 3043
rect 283 3009 330 3043
rect 168 2975 364 3009
rect 202 2941 249 2975
rect 283 2941 330 2975
rect 168 2907 364 2941
rect 202 2873 249 2907
rect 283 2873 330 2907
rect 168 2839 364 2873
rect 202 2805 249 2839
rect 283 2805 330 2839
rect 168 2771 364 2805
rect 202 2737 249 2771
rect 283 2737 330 2771
rect 168 2703 364 2737
rect 202 2669 249 2703
rect 283 2669 330 2703
rect 168 2635 364 2669
rect 202 2601 249 2635
rect 283 2601 330 2635
rect 168 2567 364 2601
rect 202 2533 249 2567
rect 283 2533 330 2567
rect 168 2499 364 2533
rect 202 2465 249 2499
rect 283 2465 330 2499
rect 168 2431 364 2465
rect 202 2397 249 2431
rect 283 2397 330 2431
rect 168 2363 364 2397
rect 202 2329 249 2363
rect 283 2329 330 2363
rect 168 2295 364 2329
rect 202 2261 249 2295
rect 283 2261 330 2295
rect 168 2227 364 2261
rect 202 2193 249 2227
rect 283 2193 330 2227
rect 168 2159 364 2193
rect 202 2125 249 2159
rect 283 2125 330 2159
rect 168 2091 364 2125
rect 202 2057 249 2091
rect 283 2057 330 2091
rect 168 2023 364 2057
rect 202 1989 249 2023
rect 283 1989 330 2023
rect 168 1955 364 1989
rect 202 1921 249 1955
rect 283 1921 330 1955
rect 168 1887 364 1921
rect 202 1853 249 1887
rect 283 1853 330 1887
rect 168 1819 364 1853
rect 202 1785 249 1819
rect 283 1785 330 1819
rect 168 1751 364 1785
rect 202 1717 249 1751
rect 283 1717 330 1751
rect 168 1683 364 1717
rect 202 1649 249 1683
rect 283 1649 330 1683
rect 168 1615 364 1649
rect 202 1581 249 1615
rect 283 1581 330 1615
rect 168 1547 364 1581
rect 202 1513 249 1547
rect 283 1513 330 1547
rect 168 1479 364 1513
rect 202 1445 249 1479
rect 283 1445 330 1479
rect 168 1411 364 1445
rect 202 1377 249 1411
rect 283 1377 330 1411
rect 168 1343 364 1377
rect 202 1309 249 1343
rect 283 1309 330 1343
rect 168 1275 364 1309
rect 202 1241 249 1275
rect 283 1241 330 1275
rect 168 1207 364 1241
rect 202 1173 249 1207
rect 283 1173 330 1207
rect 168 1139 364 1173
rect 202 1105 249 1139
rect 283 1105 330 1139
rect 168 1071 364 1105
rect 202 1037 249 1071
rect 283 1037 330 1071
rect 168 1003 364 1037
rect 202 969 249 1003
rect 283 969 330 1003
rect 168 935 364 969
rect 202 901 249 935
rect 283 901 330 935
rect 168 867 364 901
rect 202 833 249 867
rect 283 833 330 867
rect 168 799 364 833
rect 202 765 249 799
rect 283 765 330 799
rect 168 731 364 765
rect 202 697 249 731
rect 283 697 330 731
rect 168 663 364 697
rect 202 629 249 663
rect 283 629 330 663
rect 168 595 364 629
rect 202 561 249 595
rect 283 561 330 595
rect 168 527 364 561
rect 202 493 249 527
rect 283 493 330 527
rect 168 459 364 493
rect 202 425 249 459
rect 283 425 330 459
rect 168 391 364 425
rect 202 357 249 391
rect 283 357 330 391
rect 168 323 364 357
rect 202 289 249 323
rect 283 289 330 323
rect 168 255 364 289
rect 202 221 249 255
rect 283 221 330 255
rect 168 187 364 221
rect 202 153 249 187
rect 283 153 330 187
rect 168 119 364 153
rect 202 85 249 119
rect 283 85 330 119
rect 168 51 364 85
rect 202 17 249 51
rect 283 17 330 51
rect 168 -17 364 17
rect 202 -51 249 -17
rect 283 -51 330 -17
rect 168 -85 364 -51
rect 202 -119 249 -85
rect 283 -119 330 -85
rect 168 -153 364 -119
rect 202 -187 249 -153
rect 283 -187 330 -153
rect 168 -221 364 -187
rect 202 -255 249 -221
rect 283 -255 330 -221
rect 168 -289 364 -255
rect 202 -323 249 -289
rect 283 -323 330 -289
rect 168 -357 364 -323
rect 202 -391 249 -357
rect 283 -391 330 -357
rect 168 -425 364 -391
rect 202 -459 249 -425
rect 283 -459 330 -425
rect 168 -493 364 -459
rect 202 -527 249 -493
rect 283 -527 330 -493
rect 168 -561 364 -527
rect 202 -595 249 -561
rect 283 -595 330 -561
rect 168 -629 364 -595
rect 202 -663 249 -629
rect 283 -663 330 -629
rect 168 -697 364 -663
rect 202 -731 249 -697
rect 283 -731 330 -697
rect 168 -765 364 -731
rect 202 -799 249 -765
rect 283 -799 330 -765
rect 168 -833 364 -799
rect 202 -867 249 -833
rect 283 -867 330 -833
rect 168 -901 364 -867
rect 202 -935 249 -901
rect 283 -935 330 -901
rect 168 -969 364 -935
rect 202 -1003 249 -969
rect 283 -1003 330 -969
rect 168 -1037 364 -1003
rect 202 -1071 249 -1037
rect 283 -1071 330 -1037
rect 168 -1105 364 -1071
rect 202 -1139 249 -1105
rect 283 -1139 330 -1105
rect 168 -1173 364 -1139
rect 202 -1207 249 -1173
rect 283 -1207 330 -1173
rect 168 -1241 364 -1207
rect 202 -1275 249 -1241
rect 283 -1275 330 -1241
rect 168 -1309 364 -1275
rect 202 -1343 249 -1309
rect 283 -1343 330 -1309
rect 168 -1377 364 -1343
rect 202 -1411 249 -1377
rect 283 -1411 330 -1377
rect 168 -1445 364 -1411
rect 202 -1479 249 -1445
rect 283 -1479 330 -1445
rect 168 -1513 364 -1479
rect 202 -1547 249 -1513
rect 283 -1547 330 -1513
rect 168 -1581 364 -1547
rect 202 -1615 249 -1581
rect 283 -1615 330 -1581
rect 168 -1649 364 -1615
rect 202 -1683 249 -1649
rect 283 -1683 330 -1649
rect 168 -1717 364 -1683
rect 202 -1751 249 -1717
rect 283 -1751 330 -1717
rect 168 -1785 364 -1751
rect 202 -1819 249 -1785
rect 283 -1819 330 -1785
rect 168 -1853 364 -1819
rect 202 -1887 249 -1853
rect 283 -1887 330 -1853
rect 168 -1921 364 -1887
rect 202 -1955 249 -1921
rect 283 -1955 330 -1921
rect 168 -1989 364 -1955
rect 202 -2023 249 -1989
rect 283 -2023 330 -1989
rect 168 -2057 364 -2023
rect 202 -2091 249 -2057
rect 283 -2091 330 -2057
rect 168 -2125 364 -2091
rect 202 -2159 249 -2125
rect 283 -2159 330 -2125
rect 168 -2193 364 -2159
rect 202 -2227 249 -2193
rect 283 -2227 330 -2193
rect 168 -2261 364 -2227
rect 202 -2295 249 -2261
rect 283 -2295 330 -2261
rect 168 -2329 364 -2295
rect 202 -2363 249 -2329
rect 283 -2363 330 -2329
rect 168 -2397 364 -2363
rect 202 -2431 249 -2397
rect 283 -2431 330 -2397
rect 168 -2465 364 -2431
rect 202 -2499 249 -2465
rect 283 -2499 330 -2465
rect 168 -2533 364 -2499
rect 202 -2567 249 -2533
rect 283 -2567 330 -2533
rect 168 -2601 364 -2567
rect 202 -2635 249 -2601
rect 283 -2635 330 -2601
rect 168 -2669 364 -2635
rect 202 -2703 249 -2669
rect 283 -2703 330 -2669
rect 168 -2737 364 -2703
rect 202 -2771 249 -2737
rect 283 -2771 330 -2737
rect 168 -2805 364 -2771
rect 202 -2839 249 -2805
rect 283 -2839 330 -2805
rect 168 -2873 364 -2839
rect 202 -2907 249 -2873
rect 283 -2907 330 -2873
rect 168 -2941 364 -2907
rect 202 -2975 249 -2941
rect 283 -2975 330 -2941
rect 168 -3009 364 -2975
rect 202 -3043 249 -3009
rect 283 -3043 330 -3009
rect 168 -3077 364 -3043
rect 202 -3111 249 -3077
rect 283 -3111 330 -3077
rect 168 -3145 364 -3111
rect 202 -3179 249 -3145
rect 283 -3179 330 -3145
rect 168 -3213 364 -3179
rect 202 -3247 249 -3213
rect 283 -3247 330 -3213
rect 168 -3281 364 -3247
rect 202 -3315 249 -3281
rect 283 -3315 330 -3281
rect 168 -3349 364 -3315
rect 202 -3383 249 -3349
rect 283 -3383 330 -3349
rect 168 -3417 364 -3383
rect 202 -3451 249 -3417
rect 283 -3451 330 -3417
rect 168 -3485 364 -3451
rect 202 -3519 249 -3485
rect 283 -3519 330 -3485
rect 168 -3553 364 -3519
rect 202 -3587 249 -3553
rect 283 -3587 330 -3553
rect 168 -3621 364 -3587
rect 202 -3655 249 -3621
rect 283 -3655 330 -3621
rect 168 -3689 364 -3655
rect 202 -3723 249 -3689
rect 283 -3723 330 -3689
rect 168 -3757 364 -3723
rect 202 -3791 249 -3757
rect 283 -3791 330 -3757
rect 168 -3825 364 -3791
rect 202 -3859 249 -3825
rect 283 -3859 330 -3825
rect 168 -3893 364 -3859
rect 202 -3927 249 -3893
rect 283 -3927 330 -3893
rect 168 -3961 364 -3927
rect 202 -3995 249 -3961
rect 283 -3995 330 -3961
rect 168 -4029 364 -3995
rect 202 -4063 249 -4029
rect 283 -4063 330 -4029
rect 168 -4097 364 -4063
rect 202 -4131 249 -4097
rect 283 -4131 330 -4097
rect 168 -4165 364 -4131
rect 202 -4199 249 -4165
rect 283 -4199 330 -4165
rect 168 -4233 364 -4199
rect 202 -4267 249 -4233
rect 283 -4267 330 -4233
rect 168 -4301 364 -4267
rect 202 -4335 249 -4301
rect 283 -4335 330 -4301
rect 168 -4369 364 -4335
rect 202 -4403 249 -4369
rect 283 -4403 330 -4369
rect 168 -4437 364 -4403
rect 202 -4471 249 -4437
rect 283 -4471 330 -4437
rect 168 -4505 364 -4471
rect 202 -4539 249 -4505
rect 283 -4539 330 -4505
rect 168 -4573 364 -4539
rect 202 -4607 249 -4573
rect 283 -4607 330 -4573
rect 168 -4641 364 -4607
rect 202 -4675 249 -4641
rect 283 -4675 330 -4641
rect 168 -4709 364 -4675
rect 202 -4743 249 -4709
rect 283 -4743 330 -4709
rect 168 -4777 364 -4743
rect 202 -4811 249 -4777
rect 283 -4811 330 -4777
rect 168 -4845 364 -4811
rect 202 -4879 249 -4845
rect 283 -4879 330 -4845
rect 168 -4913 364 -4879
rect 202 -4947 249 -4913
rect 283 -4947 330 -4913
rect 168 -4981 364 -4947
rect -364 -5068 -168 -5015
rect 202 -5015 249 -4981
rect 283 -5015 330 -4981
rect 734 4981 781 5015
rect 815 4981 862 5015
rect 1232 5015 1330 5068
rect 700 4947 896 4981
rect 734 4913 781 4947
rect 815 4913 862 4947
rect 700 4879 896 4913
rect 734 4845 781 4879
rect 815 4845 862 4879
rect 700 4811 896 4845
rect 734 4777 781 4811
rect 815 4777 862 4811
rect 700 4743 896 4777
rect 734 4709 781 4743
rect 815 4709 862 4743
rect 700 4675 896 4709
rect 734 4641 781 4675
rect 815 4641 862 4675
rect 700 4607 896 4641
rect 734 4573 781 4607
rect 815 4573 862 4607
rect 700 4539 896 4573
rect 734 4505 781 4539
rect 815 4505 862 4539
rect 700 4471 896 4505
rect 734 4437 781 4471
rect 815 4437 862 4471
rect 700 4403 896 4437
rect 734 4369 781 4403
rect 815 4369 862 4403
rect 700 4335 896 4369
rect 734 4301 781 4335
rect 815 4301 862 4335
rect 700 4267 896 4301
rect 734 4233 781 4267
rect 815 4233 862 4267
rect 700 4199 896 4233
rect 734 4165 781 4199
rect 815 4165 862 4199
rect 700 4131 896 4165
rect 734 4097 781 4131
rect 815 4097 862 4131
rect 700 4063 896 4097
rect 734 4029 781 4063
rect 815 4029 862 4063
rect 700 3995 896 4029
rect 734 3961 781 3995
rect 815 3961 862 3995
rect 700 3927 896 3961
rect 734 3893 781 3927
rect 815 3893 862 3927
rect 700 3859 896 3893
rect 734 3825 781 3859
rect 815 3825 862 3859
rect 700 3791 896 3825
rect 734 3757 781 3791
rect 815 3757 862 3791
rect 700 3723 896 3757
rect 734 3689 781 3723
rect 815 3689 862 3723
rect 700 3655 896 3689
rect 734 3621 781 3655
rect 815 3621 862 3655
rect 700 3587 896 3621
rect 734 3553 781 3587
rect 815 3553 862 3587
rect 700 3519 896 3553
rect 734 3485 781 3519
rect 815 3485 862 3519
rect 700 3451 896 3485
rect 734 3417 781 3451
rect 815 3417 862 3451
rect 700 3383 896 3417
rect 734 3349 781 3383
rect 815 3349 862 3383
rect 700 3315 896 3349
rect 734 3281 781 3315
rect 815 3281 862 3315
rect 700 3247 896 3281
rect 734 3213 781 3247
rect 815 3213 862 3247
rect 700 3179 896 3213
rect 734 3145 781 3179
rect 815 3145 862 3179
rect 700 3111 896 3145
rect 734 3077 781 3111
rect 815 3077 862 3111
rect 700 3043 896 3077
rect 734 3009 781 3043
rect 815 3009 862 3043
rect 700 2975 896 3009
rect 734 2941 781 2975
rect 815 2941 862 2975
rect 700 2907 896 2941
rect 734 2873 781 2907
rect 815 2873 862 2907
rect 700 2839 896 2873
rect 734 2805 781 2839
rect 815 2805 862 2839
rect 700 2771 896 2805
rect 734 2737 781 2771
rect 815 2737 862 2771
rect 700 2703 896 2737
rect 734 2669 781 2703
rect 815 2669 862 2703
rect 700 2635 896 2669
rect 734 2601 781 2635
rect 815 2601 862 2635
rect 700 2567 896 2601
rect 734 2533 781 2567
rect 815 2533 862 2567
rect 700 2499 896 2533
rect 734 2465 781 2499
rect 815 2465 862 2499
rect 700 2431 896 2465
rect 734 2397 781 2431
rect 815 2397 862 2431
rect 700 2363 896 2397
rect 734 2329 781 2363
rect 815 2329 862 2363
rect 700 2295 896 2329
rect 734 2261 781 2295
rect 815 2261 862 2295
rect 700 2227 896 2261
rect 734 2193 781 2227
rect 815 2193 862 2227
rect 700 2159 896 2193
rect 734 2125 781 2159
rect 815 2125 862 2159
rect 700 2091 896 2125
rect 734 2057 781 2091
rect 815 2057 862 2091
rect 700 2023 896 2057
rect 734 1989 781 2023
rect 815 1989 862 2023
rect 700 1955 896 1989
rect 734 1921 781 1955
rect 815 1921 862 1955
rect 700 1887 896 1921
rect 734 1853 781 1887
rect 815 1853 862 1887
rect 700 1819 896 1853
rect 734 1785 781 1819
rect 815 1785 862 1819
rect 700 1751 896 1785
rect 734 1717 781 1751
rect 815 1717 862 1751
rect 700 1683 896 1717
rect 734 1649 781 1683
rect 815 1649 862 1683
rect 700 1615 896 1649
rect 734 1581 781 1615
rect 815 1581 862 1615
rect 700 1547 896 1581
rect 734 1513 781 1547
rect 815 1513 862 1547
rect 700 1479 896 1513
rect 734 1445 781 1479
rect 815 1445 862 1479
rect 700 1411 896 1445
rect 734 1377 781 1411
rect 815 1377 862 1411
rect 700 1343 896 1377
rect 734 1309 781 1343
rect 815 1309 862 1343
rect 700 1275 896 1309
rect 734 1241 781 1275
rect 815 1241 862 1275
rect 700 1207 896 1241
rect 734 1173 781 1207
rect 815 1173 862 1207
rect 700 1139 896 1173
rect 734 1105 781 1139
rect 815 1105 862 1139
rect 700 1071 896 1105
rect 734 1037 781 1071
rect 815 1037 862 1071
rect 700 1003 896 1037
rect 734 969 781 1003
rect 815 969 862 1003
rect 700 935 896 969
rect 734 901 781 935
rect 815 901 862 935
rect 700 867 896 901
rect 734 833 781 867
rect 815 833 862 867
rect 700 799 896 833
rect 734 765 781 799
rect 815 765 862 799
rect 700 731 896 765
rect 734 697 781 731
rect 815 697 862 731
rect 700 663 896 697
rect 734 629 781 663
rect 815 629 862 663
rect 700 595 896 629
rect 734 561 781 595
rect 815 561 862 595
rect 700 527 896 561
rect 734 493 781 527
rect 815 493 862 527
rect 700 459 896 493
rect 734 425 781 459
rect 815 425 862 459
rect 700 391 896 425
rect 734 357 781 391
rect 815 357 862 391
rect 700 323 896 357
rect 734 289 781 323
rect 815 289 862 323
rect 700 255 896 289
rect 734 221 781 255
rect 815 221 862 255
rect 700 187 896 221
rect 734 153 781 187
rect 815 153 862 187
rect 700 119 896 153
rect 734 85 781 119
rect 815 85 862 119
rect 700 51 896 85
rect 734 17 781 51
rect 815 17 862 51
rect 700 -17 896 17
rect 734 -51 781 -17
rect 815 -51 862 -17
rect 700 -85 896 -51
rect 734 -119 781 -85
rect 815 -119 862 -85
rect 700 -153 896 -119
rect 734 -187 781 -153
rect 815 -187 862 -153
rect 700 -221 896 -187
rect 734 -255 781 -221
rect 815 -255 862 -221
rect 700 -289 896 -255
rect 734 -323 781 -289
rect 815 -323 862 -289
rect 700 -357 896 -323
rect 734 -391 781 -357
rect 815 -391 862 -357
rect 700 -425 896 -391
rect 734 -459 781 -425
rect 815 -459 862 -425
rect 700 -493 896 -459
rect 734 -527 781 -493
rect 815 -527 862 -493
rect 700 -561 896 -527
rect 734 -595 781 -561
rect 815 -595 862 -561
rect 700 -629 896 -595
rect 734 -663 781 -629
rect 815 -663 862 -629
rect 700 -697 896 -663
rect 734 -731 781 -697
rect 815 -731 862 -697
rect 700 -765 896 -731
rect 734 -799 781 -765
rect 815 -799 862 -765
rect 700 -833 896 -799
rect 734 -867 781 -833
rect 815 -867 862 -833
rect 700 -901 896 -867
rect 734 -935 781 -901
rect 815 -935 862 -901
rect 700 -969 896 -935
rect 734 -1003 781 -969
rect 815 -1003 862 -969
rect 700 -1037 896 -1003
rect 734 -1071 781 -1037
rect 815 -1071 862 -1037
rect 700 -1105 896 -1071
rect 734 -1139 781 -1105
rect 815 -1139 862 -1105
rect 700 -1173 896 -1139
rect 734 -1207 781 -1173
rect 815 -1207 862 -1173
rect 700 -1241 896 -1207
rect 734 -1275 781 -1241
rect 815 -1275 862 -1241
rect 700 -1309 896 -1275
rect 734 -1343 781 -1309
rect 815 -1343 862 -1309
rect 700 -1377 896 -1343
rect 734 -1411 781 -1377
rect 815 -1411 862 -1377
rect 700 -1445 896 -1411
rect 734 -1479 781 -1445
rect 815 -1479 862 -1445
rect 700 -1513 896 -1479
rect 734 -1547 781 -1513
rect 815 -1547 862 -1513
rect 700 -1581 896 -1547
rect 734 -1615 781 -1581
rect 815 -1615 862 -1581
rect 700 -1649 896 -1615
rect 734 -1683 781 -1649
rect 815 -1683 862 -1649
rect 700 -1717 896 -1683
rect 734 -1751 781 -1717
rect 815 -1751 862 -1717
rect 700 -1785 896 -1751
rect 734 -1819 781 -1785
rect 815 -1819 862 -1785
rect 700 -1853 896 -1819
rect 734 -1887 781 -1853
rect 815 -1887 862 -1853
rect 700 -1921 896 -1887
rect 734 -1955 781 -1921
rect 815 -1955 862 -1921
rect 700 -1989 896 -1955
rect 734 -2023 781 -1989
rect 815 -2023 862 -1989
rect 700 -2057 896 -2023
rect 734 -2091 781 -2057
rect 815 -2091 862 -2057
rect 700 -2125 896 -2091
rect 734 -2159 781 -2125
rect 815 -2159 862 -2125
rect 700 -2193 896 -2159
rect 734 -2227 781 -2193
rect 815 -2227 862 -2193
rect 700 -2261 896 -2227
rect 734 -2295 781 -2261
rect 815 -2295 862 -2261
rect 700 -2329 896 -2295
rect 734 -2363 781 -2329
rect 815 -2363 862 -2329
rect 700 -2397 896 -2363
rect 734 -2431 781 -2397
rect 815 -2431 862 -2397
rect 700 -2465 896 -2431
rect 734 -2499 781 -2465
rect 815 -2499 862 -2465
rect 700 -2533 896 -2499
rect 734 -2567 781 -2533
rect 815 -2567 862 -2533
rect 700 -2601 896 -2567
rect 734 -2635 781 -2601
rect 815 -2635 862 -2601
rect 700 -2669 896 -2635
rect 734 -2703 781 -2669
rect 815 -2703 862 -2669
rect 700 -2737 896 -2703
rect 734 -2771 781 -2737
rect 815 -2771 862 -2737
rect 700 -2805 896 -2771
rect 734 -2839 781 -2805
rect 815 -2839 862 -2805
rect 700 -2873 896 -2839
rect 734 -2907 781 -2873
rect 815 -2907 862 -2873
rect 700 -2941 896 -2907
rect 734 -2975 781 -2941
rect 815 -2975 862 -2941
rect 700 -3009 896 -2975
rect 734 -3043 781 -3009
rect 815 -3043 862 -3009
rect 700 -3077 896 -3043
rect 734 -3111 781 -3077
rect 815 -3111 862 -3077
rect 700 -3145 896 -3111
rect 734 -3179 781 -3145
rect 815 -3179 862 -3145
rect 700 -3213 896 -3179
rect 734 -3247 781 -3213
rect 815 -3247 862 -3213
rect 700 -3281 896 -3247
rect 734 -3315 781 -3281
rect 815 -3315 862 -3281
rect 700 -3349 896 -3315
rect 734 -3383 781 -3349
rect 815 -3383 862 -3349
rect 700 -3417 896 -3383
rect 734 -3451 781 -3417
rect 815 -3451 862 -3417
rect 700 -3485 896 -3451
rect 734 -3519 781 -3485
rect 815 -3519 862 -3485
rect 700 -3553 896 -3519
rect 734 -3587 781 -3553
rect 815 -3587 862 -3553
rect 700 -3621 896 -3587
rect 734 -3655 781 -3621
rect 815 -3655 862 -3621
rect 700 -3689 896 -3655
rect 734 -3723 781 -3689
rect 815 -3723 862 -3689
rect 700 -3757 896 -3723
rect 734 -3791 781 -3757
rect 815 -3791 862 -3757
rect 700 -3825 896 -3791
rect 734 -3859 781 -3825
rect 815 -3859 862 -3825
rect 700 -3893 896 -3859
rect 734 -3927 781 -3893
rect 815 -3927 862 -3893
rect 700 -3961 896 -3927
rect 734 -3995 781 -3961
rect 815 -3995 862 -3961
rect 700 -4029 896 -3995
rect 734 -4063 781 -4029
rect 815 -4063 862 -4029
rect 700 -4097 896 -4063
rect 734 -4131 781 -4097
rect 815 -4131 862 -4097
rect 700 -4165 896 -4131
rect 734 -4199 781 -4165
rect 815 -4199 862 -4165
rect 700 -4233 896 -4199
rect 734 -4267 781 -4233
rect 815 -4267 862 -4233
rect 700 -4301 896 -4267
rect 734 -4335 781 -4301
rect 815 -4335 862 -4301
rect 700 -4369 896 -4335
rect 734 -4403 781 -4369
rect 815 -4403 862 -4369
rect 700 -4437 896 -4403
rect 734 -4471 781 -4437
rect 815 -4471 862 -4437
rect 700 -4505 896 -4471
rect 734 -4539 781 -4505
rect 815 -4539 862 -4505
rect 700 -4573 896 -4539
rect 734 -4607 781 -4573
rect 815 -4607 862 -4573
rect 700 -4641 896 -4607
rect 734 -4675 781 -4641
rect 815 -4675 862 -4641
rect 700 -4709 896 -4675
rect 734 -4743 781 -4709
rect 815 -4743 862 -4709
rect 700 -4777 896 -4743
rect 734 -4811 781 -4777
rect 815 -4811 862 -4777
rect 700 -4845 896 -4811
rect 734 -4879 781 -4845
rect 815 -4879 862 -4845
rect 700 -4913 896 -4879
rect 734 -4947 781 -4913
rect 815 -4947 862 -4913
rect 700 -4981 896 -4947
rect 168 -5068 364 -5015
rect 734 -5015 781 -4981
rect 815 -5015 862 -4981
rect 1266 4981 1330 5015
rect 1232 4947 1330 4981
rect 1266 4913 1330 4947
rect 1232 4879 1330 4913
rect 1266 4845 1330 4879
rect 1232 4811 1330 4845
rect 1266 4777 1330 4811
rect 1232 4743 1330 4777
rect 1266 4709 1330 4743
rect 1232 4675 1330 4709
rect 1266 4641 1330 4675
rect 1232 4607 1330 4641
rect 1266 4573 1330 4607
rect 1232 4539 1330 4573
rect 1266 4505 1330 4539
rect 1232 4471 1330 4505
rect 1266 4437 1330 4471
rect 1232 4403 1330 4437
rect 1266 4369 1330 4403
rect 1232 4335 1330 4369
rect 1266 4301 1330 4335
rect 1232 4267 1330 4301
rect 1266 4233 1330 4267
rect 1232 4199 1330 4233
rect 1266 4165 1330 4199
rect 1232 4131 1330 4165
rect 1266 4097 1330 4131
rect 1232 4063 1330 4097
rect 1266 4029 1330 4063
rect 1232 3995 1330 4029
rect 1266 3961 1330 3995
rect 1232 3927 1330 3961
rect 1266 3893 1330 3927
rect 1232 3859 1330 3893
rect 1266 3825 1330 3859
rect 1232 3791 1330 3825
rect 1266 3757 1330 3791
rect 1232 3723 1330 3757
rect 1266 3689 1330 3723
rect 1232 3655 1330 3689
rect 1266 3621 1330 3655
rect 1232 3587 1330 3621
rect 1266 3553 1330 3587
rect 1232 3519 1330 3553
rect 1266 3485 1330 3519
rect 1232 3451 1330 3485
rect 1266 3417 1330 3451
rect 1232 3383 1330 3417
rect 1266 3349 1330 3383
rect 1232 3315 1330 3349
rect 1266 3281 1330 3315
rect 1232 3247 1330 3281
rect 1266 3213 1330 3247
rect 1232 3179 1330 3213
rect 1266 3145 1330 3179
rect 1232 3111 1330 3145
rect 1266 3077 1330 3111
rect 1232 3043 1330 3077
rect 1266 3009 1330 3043
rect 1232 2975 1330 3009
rect 1266 2941 1330 2975
rect 1232 2907 1330 2941
rect 1266 2873 1330 2907
rect 1232 2839 1330 2873
rect 1266 2805 1330 2839
rect 1232 2771 1330 2805
rect 1266 2737 1330 2771
rect 1232 2703 1330 2737
rect 1266 2669 1330 2703
rect 1232 2635 1330 2669
rect 1266 2601 1330 2635
rect 1232 2567 1330 2601
rect 1266 2533 1330 2567
rect 1232 2499 1330 2533
rect 1266 2465 1330 2499
rect 1232 2431 1330 2465
rect 1266 2397 1330 2431
rect 1232 2363 1330 2397
rect 1266 2329 1330 2363
rect 1232 2295 1330 2329
rect 1266 2261 1330 2295
rect 1232 2227 1330 2261
rect 1266 2193 1330 2227
rect 1232 2159 1330 2193
rect 1266 2125 1330 2159
rect 1232 2091 1330 2125
rect 1266 2057 1330 2091
rect 1232 2023 1330 2057
rect 1266 1989 1330 2023
rect 1232 1955 1330 1989
rect 1266 1921 1330 1955
rect 1232 1887 1330 1921
rect 1266 1853 1330 1887
rect 1232 1819 1330 1853
rect 1266 1785 1330 1819
rect 1232 1751 1330 1785
rect 1266 1717 1330 1751
rect 1232 1683 1330 1717
rect 1266 1649 1330 1683
rect 1232 1615 1330 1649
rect 1266 1581 1330 1615
rect 1232 1547 1330 1581
rect 1266 1513 1330 1547
rect 1232 1479 1330 1513
rect 1266 1445 1330 1479
rect 1232 1411 1330 1445
rect 1266 1377 1330 1411
rect 1232 1343 1330 1377
rect 1266 1309 1330 1343
rect 1232 1275 1330 1309
rect 1266 1241 1330 1275
rect 1232 1207 1330 1241
rect 1266 1173 1330 1207
rect 1232 1139 1330 1173
rect 1266 1105 1330 1139
rect 1232 1071 1330 1105
rect 1266 1037 1330 1071
rect 1232 1003 1330 1037
rect 1266 969 1330 1003
rect 1232 935 1330 969
rect 1266 901 1330 935
rect 1232 867 1330 901
rect 1266 833 1330 867
rect 1232 799 1330 833
rect 1266 765 1330 799
rect 1232 731 1330 765
rect 1266 697 1330 731
rect 1232 663 1330 697
rect 1266 629 1330 663
rect 1232 595 1330 629
rect 1266 561 1330 595
rect 1232 527 1330 561
rect 1266 493 1330 527
rect 1232 459 1330 493
rect 1266 425 1330 459
rect 1232 391 1330 425
rect 1266 357 1330 391
rect 1232 323 1330 357
rect 1266 289 1330 323
rect 1232 255 1330 289
rect 1266 221 1330 255
rect 1232 187 1330 221
rect 1266 153 1330 187
rect 1232 119 1330 153
rect 1266 85 1330 119
rect 1232 51 1330 85
rect 1266 17 1330 51
rect 1232 -17 1330 17
rect 1266 -51 1330 -17
rect 1232 -85 1330 -51
rect 1266 -119 1330 -85
rect 1232 -153 1330 -119
rect 1266 -187 1330 -153
rect 1232 -221 1330 -187
rect 1266 -255 1330 -221
rect 1232 -289 1330 -255
rect 1266 -323 1330 -289
rect 1232 -357 1330 -323
rect 1266 -391 1330 -357
rect 1232 -425 1330 -391
rect 1266 -459 1330 -425
rect 1232 -493 1330 -459
rect 1266 -527 1330 -493
rect 1232 -561 1330 -527
rect 1266 -595 1330 -561
rect 1232 -629 1330 -595
rect 1266 -663 1330 -629
rect 1232 -697 1330 -663
rect 1266 -731 1330 -697
rect 1232 -765 1330 -731
rect 1266 -799 1330 -765
rect 1232 -833 1330 -799
rect 1266 -867 1330 -833
rect 1232 -901 1330 -867
rect 1266 -935 1330 -901
rect 1232 -969 1330 -935
rect 1266 -1003 1330 -969
rect 1232 -1037 1330 -1003
rect 1266 -1071 1330 -1037
rect 1232 -1105 1330 -1071
rect 1266 -1139 1330 -1105
rect 1232 -1173 1330 -1139
rect 1266 -1207 1330 -1173
rect 1232 -1241 1330 -1207
rect 1266 -1275 1330 -1241
rect 1232 -1309 1330 -1275
rect 1266 -1343 1330 -1309
rect 1232 -1377 1330 -1343
rect 1266 -1411 1330 -1377
rect 1232 -1445 1330 -1411
rect 1266 -1479 1330 -1445
rect 1232 -1513 1330 -1479
rect 1266 -1547 1330 -1513
rect 1232 -1581 1330 -1547
rect 1266 -1615 1330 -1581
rect 1232 -1649 1330 -1615
rect 1266 -1683 1330 -1649
rect 1232 -1717 1330 -1683
rect 1266 -1751 1330 -1717
rect 1232 -1785 1330 -1751
rect 1266 -1819 1330 -1785
rect 1232 -1853 1330 -1819
rect 1266 -1887 1330 -1853
rect 1232 -1921 1330 -1887
rect 1266 -1955 1330 -1921
rect 1232 -1989 1330 -1955
rect 1266 -2023 1330 -1989
rect 1232 -2057 1330 -2023
rect 1266 -2091 1330 -2057
rect 1232 -2125 1330 -2091
rect 1266 -2159 1330 -2125
rect 1232 -2193 1330 -2159
rect 1266 -2227 1330 -2193
rect 1232 -2261 1330 -2227
rect 1266 -2295 1330 -2261
rect 1232 -2329 1330 -2295
rect 1266 -2363 1330 -2329
rect 1232 -2397 1330 -2363
rect 1266 -2431 1330 -2397
rect 1232 -2465 1330 -2431
rect 1266 -2499 1330 -2465
rect 1232 -2533 1330 -2499
rect 1266 -2567 1330 -2533
rect 1232 -2601 1330 -2567
rect 1266 -2635 1330 -2601
rect 1232 -2669 1330 -2635
rect 1266 -2703 1330 -2669
rect 1232 -2737 1330 -2703
rect 1266 -2771 1330 -2737
rect 1232 -2805 1330 -2771
rect 1266 -2839 1330 -2805
rect 1232 -2873 1330 -2839
rect 1266 -2907 1330 -2873
rect 1232 -2941 1330 -2907
rect 1266 -2975 1330 -2941
rect 1232 -3009 1330 -2975
rect 1266 -3043 1330 -3009
rect 1232 -3077 1330 -3043
rect 1266 -3111 1330 -3077
rect 1232 -3145 1330 -3111
rect 1266 -3179 1330 -3145
rect 1232 -3213 1330 -3179
rect 1266 -3247 1330 -3213
rect 1232 -3281 1330 -3247
rect 1266 -3315 1330 -3281
rect 1232 -3349 1330 -3315
rect 1266 -3383 1330 -3349
rect 1232 -3417 1330 -3383
rect 1266 -3451 1330 -3417
rect 1232 -3485 1330 -3451
rect 1266 -3519 1330 -3485
rect 1232 -3553 1330 -3519
rect 1266 -3587 1330 -3553
rect 1232 -3621 1330 -3587
rect 1266 -3655 1330 -3621
rect 1232 -3689 1330 -3655
rect 1266 -3723 1330 -3689
rect 1232 -3757 1330 -3723
rect 1266 -3791 1330 -3757
rect 1232 -3825 1330 -3791
rect 1266 -3859 1330 -3825
rect 1232 -3893 1330 -3859
rect 1266 -3927 1330 -3893
rect 1232 -3961 1330 -3927
rect 1266 -3995 1330 -3961
rect 1232 -4029 1330 -3995
rect 1266 -4063 1330 -4029
rect 1232 -4097 1330 -4063
rect 1266 -4131 1330 -4097
rect 1232 -4165 1330 -4131
rect 1266 -4199 1330 -4165
rect 1232 -4233 1330 -4199
rect 1266 -4267 1330 -4233
rect 1232 -4301 1330 -4267
rect 1266 -4335 1330 -4301
rect 1232 -4369 1330 -4335
rect 1266 -4403 1330 -4369
rect 1232 -4437 1330 -4403
rect 1266 -4471 1330 -4437
rect 1232 -4505 1330 -4471
rect 1266 -4539 1330 -4505
rect 1232 -4573 1330 -4539
rect 1266 -4607 1330 -4573
rect 1232 -4641 1330 -4607
rect 1266 -4675 1330 -4641
rect 1232 -4709 1330 -4675
rect 1266 -4743 1330 -4709
rect 1232 -4777 1330 -4743
rect 1266 -4811 1330 -4777
rect 1232 -4845 1330 -4811
rect 1266 -4879 1330 -4845
rect 1232 -4913 1330 -4879
rect 1266 -4947 1330 -4913
rect 1232 -4981 1330 -4947
rect 700 -5068 896 -5015
rect 1266 -5015 1330 -4981
rect 1232 -5068 1330 -5015
rect -1330 -5102 -1183 -5068
rect -1149 -5102 -1115 -5068
rect -1081 -5102 -1047 -5068
rect -1013 -5102 -979 -5068
rect -945 -5102 -651 -5068
rect -617 -5102 -583 -5068
rect -549 -5102 -515 -5068
rect -481 -5102 -447 -5068
rect -413 -5102 -119 -5068
rect -85 -5102 -51 -5068
rect -17 -5102 17 -5068
rect 51 -5102 85 -5068
rect 119 -5102 413 -5068
rect 447 -5102 481 -5068
rect 515 -5102 549 -5068
rect 583 -5102 617 -5068
rect 651 -5102 945 -5068
rect 979 -5102 1013 -5068
rect 1047 -5102 1081 -5068
rect 1115 -5102 1149 -5068
rect 1183 -5102 1330 -5068
<< mvpsubdiffcont >>
rect -1411 5356 1411 5730
rect -1926 -5219 -1552 5219
rect 1552 -5219 1926 5219
rect -1411 -5730 1411 -5356
<< mvnsubdiffcont >>
rect -1183 5068 -1149 5102
rect -1115 5068 -1081 5102
rect -1047 5068 -1013 5102
rect -979 5068 -945 5102
rect -651 5068 -617 5102
rect -583 5068 -549 5102
rect -515 5068 -481 5102
rect -447 5068 -413 5102
rect -119 5068 -85 5102
rect -51 5068 -17 5102
rect 17 5068 51 5102
rect 85 5068 119 5102
rect 413 5068 447 5102
rect 481 5068 515 5102
rect 549 5068 583 5102
rect 617 5068 651 5102
rect 945 5068 979 5102
rect 1013 5068 1047 5102
rect 1081 5068 1115 5102
rect 1149 5068 1183 5102
rect -1266 4981 -1232 5015
rect -1266 4913 -1232 4947
rect -1266 4845 -1232 4879
rect -1266 4777 -1232 4811
rect -1266 4709 -1232 4743
rect -1266 4641 -1232 4675
rect -1266 4573 -1232 4607
rect -1266 4505 -1232 4539
rect -1266 4437 -1232 4471
rect -1266 4369 -1232 4403
rect -1266 4301 -1232 4335
rect -1266 4233 -1232 4267
rect -1266 4165 -1232 4199
rect -1266 4097 -1232 4131
rect -1266 4029 -1232 4063
rect -1266 3961 -1232 3995
rect -1266 3893 -1232 3927
rect -1266 3825 -1232 3859
rect -1266 3757 -1232 3791
rect -1266 3689 -1232 3723
rect -1266 3621 -1232 3655
rect -1266 3553 -1232 3587
rect -1266 3485 -1232 3519
rect -1266 3417 -1232 3451
rect -1266 3349 -1232 3383
rect -1266 3281 -1232 3315
rect -1266 3213 -1232 3247
rect -1266 3145 -1232 3179
rect -1266 3077 -1232 3111
rect -1266 3009 -1232 3043
rect -1266 2941 -1232 2975
rect -1266 2873 -1232 2907
rect -1266 2805 -1232 2839
rect -1266 2737 -1232 2771
rect -1266 2669 -1232 2703
rect -1266 2601 -1232 2635
rect -1266 2533 -1232 2567
rect -1266 2465 -1232 2499
rect -1266 2397 -1232 2431
rect -1266 2329 -1232 2363
rect -1266 2261 -1232 2295
rect -1266 2193 -1232 2227
rect -1266 2125 -1232 2159
rect -1266 2057 -1232 2091
rect -1266 1989 -1232 2023
rect -1266 1921 -1232 1955
rect -1266 1853 -1232 1887
rect -1266 1785 -1232 1819
rect -1266 1717 -1232 1751
rect -1266 1649 -1232 1683
rect -1266 1581 -1232 1615
rect -1266 1513 -1232 1547
rect -1266 1445 -1232 1479
rect -1266 1377 -1232 1411
rect -1266 1309 -1232 1343
rect -1266 1241 -1232 1275
rect -1266 1173 -1232 1207
rect -1266 1105 -1232 1139
rect -1266 1037 -1232 1071
rect -1266 969 -1232 1003
rect -1266 901 -1232 935
rect -1266 833 -1232 867
rect -1266 765 -1232 799
rect -1266 697 -1232 731
rect -1266 629 -1232 663
rect -1266 561 -1232 595
rect -1266 493 -1232 527
rect -1266 425 -1232 459
rect -1266 357 -1232 391
rect -1266 289 -1232 323
rect -1266 221 -1232 255
rect -1266 153 -1232 187
rect -1266 85 -1232 119
rect -1266 17 -1232 51
rect -1266 -51 -1232 -17
rect -1266 -119 -1232 -85
rect -1266 -187 -1232 -153
rect -1266 -255 -1232 -221
rect -1266 -323 -1232 -289
rect -1266 -391 -1232 -357
rect -1266 -459 -1232 -425
rect -1266 -527 -1232 -493
rect -1266 -595 -1232 -561
rect -1266 -663 -1232 -629
rect -1266 -731 -1232 -697
rect -1266 -799 -1232 -765
rect -1266 -867 -1232 -833
rect -1266 -935 -1232 -901
rect -1266 -1003 -1232 -969
rect -1266 -1071 -1232 -1037
rect -1266 -1139 -1232 -1105
rect -1266 -1207 -1232 -1173
rect -1266 -1275 -1232 -1241
rect -1266 -1343 -1232 -1309
rect -1266 -1411 -1232 -1377
rect -1266 -1479 -1232 -1445
rect -1266 -1547 -1232 -1513
rect -1266 -1615 -1232 -1581
rect -1266 -1683 -1232 -1649
rect -1266 -1751 -1232 -1717
rect -1266 -1819 -1232 -1785
rect -1266 -1887 -1232 -1853
rect -1266 -1955 -1232 -1921
rect -1266 -2023 -1232 -1989
rect -1266 -2091 -1232 -2057
rect -1266 -2159 -1232 -2125
rect -1266 -2227 -1232 -2193
rect -1266 -2295 -1232 -2261
rect -1266 -2363 -1232 -2329
rect -1266 -2431 -1232 -2397
rect -1266 -2499 -1232 -2465
rect -1266 -2567 -1232 -2533
rect -1266 -2635 -1232 -2601
rect -1266 -2703 -1232 -2669
rect -1266 -2771 -1232 -2737
rect -1266 -2839 -1232 -2805
rect -1266 -2907 -1232 -2873
rect -1266 -2975 -1232 -2941
rect -1266 -3043 -1232 -3009
rect -1266 -3111 -1232 -3077
rect -1266 -3179 -1232 -3145
rect -1266 -3247 -1232 -3213
rect -1266 -3315 -1232 -3281
rect -1266 -3383 -1232 -3349
rect -1266 -3451 -1232 -3417
rect -1266 -3519 -1232 -3485
rect -1266 -3587 -1232 -3553
rect -1266 -3655 -1232 -3621
rect -1266 -3723 -1232 -3689
rect -1266 -3791 -1232 -3757
rect -1266 -3859 -1232 -3825
rect -1266 -3927 -1232 -3893
rect -1266 -3995 -1232 -3961
rect -1266 -4063 -1232 -4029
rect -1266 -4131 -1232 -4097
rect -1266 -4199 -1232 -4165
rect -1266 -4267 -1232 -4233
rect -1266 -4335 -1232 -4301
rect -1266 -4403 -1232 -4369
rect -1266 -4471 -1232 -4437
rect -1266 -4539 -1232 -4505
rect -1266 -4607 -1232 -4573
rect -1266 -4675 -1232 -4641
rect -1266 -4743 -1232 -4709
rect -1266 -4811 -1232 -4777
rect -1266 -4879 -1232 -4845
rect -1266 -4947 -1232 -4913
rect -1266 -5015 -1232 -4981
rect -896 4981 -862 5015
rect -815 4981 -781 5015
rect -734 4981 -700 5015
rect -896 4913 -862 4947
rect -815 4913 -781 4947
rect -734 4913 -700 4947
rect -896 4845 -862 4879
rect -815 4845 -781 4879
rect -734 4845 -700 4879
rect -896 4777 -862 4811
rect -815 4777 -781 4811
rect -734 4777 -700 4811
rect -896 4709 -862 4743
rect -815 4709 -781 4743
rect -734 4709 -700 4743
rect -896 4641 -862 4675
rect -815 4641 -781 4675
rect -734 4641 -700 4675
rect -896 4573 -862 4607
rect -815 4573 -781 4607
rect -734 4573 -700 4607
rect -896 4505 -862 4539
rect -815 4505 -781 4539
rect -734 4505 -700 4539
rect -896 4437 -862 4471
rect -815 4437 -781 4471
rect -734 4437 -700 4471
rect -896 4369 -862 4403
rect -815 4369 -781 4403
rect -734 4369 -700 4403
rect -896 4301 -862 4335
rect -815 4301 -781 4335
rect -734 4301 -700 4335
rect -896 4233 -862 4267
rect -815 4233 -781 4267
rect -734 4233 -700 4267
rect -896 4165 -862 4199
rect -815 4165 -781 4199
rect -734 4165 -700 4199
rect -896 4097 -862 4131
rect -815 4097 -781 4131
rect -734 4097 -700 4131
rect -896 4029 -862 4063
rect -815 4029 -781 4063
rect -734 4029 -700 4063
rect -896 3961 -862 3995
rect -815 3961 -781 3995
rect -734 3961 -700 3995
rect -896 3893 -862 3927
rect -815 3893 -781 3927
rect -734 3893 -700 3927
rect -896 3825 -862 3859
rect -815 3825 -781 3859
rect -734 3825 -700 3859
rect -896 3757 -862 3791
rect -815 3757 -781 3791
rect -734 3757 -700 3791
rect -896 3689 -862 3723
rect -815 3689 -781 3723
rect -734 3689 -700 3723
rect -896 3621 -862 3655
rect -815 3621 -781 3655
rect -734 3621 -700 3655
rect -896 3553 -862 3587
rect -815 3553 -781 3587
rect -734 3553 -700 3587
rect -896 3485 -862 3519
rect -815 3485 -781 3519
rect -734 3485 -700 3519
rect -896 3417 -862 3451
rect -815 3417 -781 3451
rect -734 3417 -700 3451
rect -896 3349 -862 3383
rect -815 3349 -781 3383
rect -734 3349 -700 3383
rect -896 3281 -862 3315
rect -815 3281 -781 3315
rect -734 3281 -700 3315
rect -896 3213 -862 3247
rect -815 3213 -781 3247
rect -734 3213 -700 3247
rect -896 3145 -862 3179
rect -815 3145 -781 3179
rect -734 3145 -700 3179
rect -896 3077 -862 3111
rect -815 3077 -781 3111
rect -734 3077 -700 3111
rect -896 3009 -862 3043
rect -815 3009 -781 3043
rect -734 3009 -700 3043
rect -896 2941 -862 2975
rect -815 2941 -781 2975
rect -734 2941 -700 2975
rect -896 2873 -862 2907
rect -815 2873 -781 2907
rect -734 2873 -700 2907
rect -896 2805 -862 2839
rect -815 2805 -781 2839
rect -734 2805 -700 2839
rect -896 2737 -862 2771
rect -815 2737 -781 2771
rect -734 2737 -700 2771
rect -896 2669 -862 2703
rect -815 2669 -781 2703
rect -734 2669 -700 2703
rect -896 2601 -862 2635
rect -815 2601 -781 2635
rect -734 2601 -700 2635
rect -896 2533 -862 2567
rect -815 2533 -781 2567
rect -734 2533 -700 2567
rect -896 2465 -862 2499
rect -815 2465 -781 2499
rect -734 2465 -700 2499
rect -896 2397 -862 2431
rect -815 2397 -781 2431
rect -734 2397 -700 2431
rect -896 2329 -862 2363
rect -815 2329 -781 2363
rect -734 2329 -700 2363
rect -896 2261 -862 2295
rect -815 2261 -781 2295
rect -734 2261 -700 2295
rect -896 2193 -862 2227
rect -815 2193 -781 2227
rect -734 2193 -700 2227
rect -896 2125 -862 2159
rect -815 2125 -781 2159
rect -734 2125 -700 2159
rect -896 2057 -862 2091
rect -815 2057 -781 2091
rect -734 2057 -700 2091
rect -896 1989 -862 2023
rect -815 1989 -781 2023
rect -734 1989 -700 2023
rect -896 1921 -862 1955
rect -815 1921 -781 1955
rect -734 1921 -700 1955
rect -896 1853 -862 1887
rect -815 1853 -781 1887
rect -734 1853 -700 1887
rect -896 1785 -862 1819
rect -815 1785 -781 1819
rect -734 1785 -700 1819
rect -896 1717 -862 1751
rect -815 1717 -781 1751
rect -734 1717 -700 1751
rect -896 1649 -862 1683
rect -815 1649 -781 1683
rect -734 1649 -700 1683
rect -896 1581 -862 1615
rect -815 1581 -781 1615
rect -734 1581 -700 1615
rect -896 1513 -862 1547
rect -815 1513 -781 1547
rect -734 1513 -700 1547
rect -896 1445 -862 1479
rect -815 1445 -781 1479
rect -734 1445 -700 1479
rect -896 1377 -862 1411
rect -815 1377 -781 1411
rect -734 1377 -700 1411
rect -896 1309 -862 1343
rect -815 1309 -781 1343
rect -734 1309 -700 1343
rect -896 1241 -862 1275
rect -815 1241 -781 1275
rect -734 1241 -700 1275
rect -896 1173 -862 1207
rect -815 1173 -781 1207
rect -734 1173 -700 1207
rect -896 1105 -862 1139
rect -815 1105 -781 1139
rect -734 1105 -700 1139
rect -896 1037 -862 1071
rect -815 1037 -781 1071
rect -734 1037 -700 1071
rect -896 969 -862 1003
rect -815 969 -781 1003
rect -734 969 -700 1003
rect -896 901 -862 935
rect -815 901 -781 935
rect -734 901 -700 935
rect -896 833 -862 867
rect -815 833 -781 867
rect -734 833 -700 867
rect -896 765 -862 799
rect -815 765 -781 799
rect -734 765 -700 799
rect -896 697 -862 731
rect -815 697 -781 731
rect -734 697 -700 731
rect -896 629 -862 663
rect -815 629 -781 663
rect -734 629 -700 663
rect -896 561 -862 595
rect -815 561 -781 595
rect -734 561 -700 595
rect -896 493 -862 527
rect -815 493 -781 527
rect -734 493 -700 527
rect -896 425 -862 459
rect -815 425 -781 459
rect -734 425 -700 459
rect -896 357 -862 391
rect -815 357 -781 391
rect -734 357 -700 391
rect -896 289 -862 323
rect -815 289 -781 323
rect -734 289 -700 323
rect -896 221 -862 255
rect -815 221 -781 255
rect -734 221 -700 255
rect -896 153 -862 187
rect -815 153 -781 187
rect -734 153 -700 187
rect -896 85 -862 119
rect -815 85 -781 119
rect -734 85 -700 119
rect -896 17 -862 51
rect -815 17 -781 51
rect -734 17 -700 51
rect -896 -51 -862 -17
rect -815 -51 -781 -17
rect -734 -51 -700 -17
rect -896 -119 -862 -85
rect -815 -119 -781 -85
rect -734 -119 -700 -85
rect -896 -187 -862 -153
rect -815 -187 -781 -153
rect -734 -187 -700 -153
rect -896 -255 -862 -221
rect -815 -255 -781 -221
rect -734 -255 -700 -221
rect -896 -323 -862 -289
rect -815 -323 -781 -289
rect -734 -323 -700 -289
rect -896 -391 -862 -357
rect -815 -391 -781 -357
rect -734 -391 -700 -357
rect -896 -459 -862 -425
rect -815 -459 -781 -425
rect -734 -459 -700 -425
rect -896 -527 -862 -493
rect -815 -527 -781 -493
rect -734 -527 -700 -493
rect -896 -595 -862 -561
rect -815 -595 -781 -561
rect -734 -595 -700 -561
rect -896 -663 -862 -629
rect -815 -663 -781 -629
rect -734 -663 -700 -629
rect -896 -731 -862 -697
rect -815 -731 -781 -697
rect -734 -731 -700 -697
rect -896 -799 -862 -765
rect -815 -799 -781 -765
rect -734 -799 -700 -765
rect -896 -867 -862 -833
rect -815 -867 -781 -833
rect -734 -867 -700 -833
rect -896 -935 -862 -901
rect -815 -935 -781 -901
rect -734 -935 -700 -901
rect -896 -1003 -862 -969
rect -815 -1003 -781 -969
rect -734 -1003 -700 -969
rect -896 -1071 -862 -1037
rect -815 -1071 -781 -1037
rect -734 -1071 -700 -1037
rect -896 -1139 -862 -1105
rect -815 -1139 -781 -1105
rect -734 -1139 -700 -1105
rect -896 -1207 -862 -1173
rect -815 -1207 -781 -1173
rect -734 -1207 -700 -1173
rect -896 -1275 -862 -1241
rect -815 -1275 -781 -1241
rect -734 -1275 -700 -1241
rect -896 -1343 -862 -1309
rect -815 -1343 -781 -1309
rect -734 -1343 -700 -1309
rect -896 -1411 -862 -1377
rect -815 -1411 -781 -1377
rect -734 -1411 -700 -1377
rect -896 -1479 -862 -1445
rect -815 -1479 -781 -1445
rect -734 -1479 -700 -1445
rect -896 -1547 -862 -1513
rect -815 -1547 -781 -1513
rect -734 -1547 -700 -1513
rect -896 -1615 -862 -1581
rect -815 -1615 -781 -1581
rect -734 -1615 -700 -1581
rect -896 -1683 -862 -1649
rect -815 -1683 -781 -1649
rect -734 -1683 -700 -1649
rect -896 -1751 -862 -1717
rect -815 -1751 -781 -1717
rect -734 -1751 -700 -1717
rect -896 -1819 -862 -1785
rect -815 -1819 -781 -1785
rect -734 -1819 -700 -1785
rect -896 -1887 -862 -1853
rect -815 -1887 -781 -1853
rect -734 -1887 -700 -1853
rect -896 -1955 -862 -1921
rect -815 -1955 -781 -1921
rect -734 -1955 -700 -1921
rect -896 -2023 -862 -1989
rect -815 -2023 -781 -1989
rect -734 -2023 -700 -1989
rect -896 -2091 -862 -2057
rect -815 -2091 -781 -2057
rect -734 -2091 -700 -2057
rect -896 -2159 -862 -2125
rect -815 -2159 -781 -2125
rect -734 -2159 -700 -2125
rect -896 -2227 -862 -2193
rect -815 -2227 -781 -2193
rect -734 -2227 -700 -2193
rect -896 -2295 -862 -2261
rect -815 -2295 -781 -2261
rect -734 -2295 -700 -2261
rect -896 -2363 -862 -2329
rect -815 -2363 -781 -2329
rect -734 -2363 -700 -2329
rect -896 -2431 -862 -2397
rect -815 -2431 -781 -2397
rect -734 -2431 -700 -2397
rect -896 -2499 -862 -2465
rect -815 -2499 -781 -2465
rect -734 -2499 -700 -2465
rect -896 -2567 -862 -2533
rect -815 -2567 -781 -2533
rect -734 -2567 -700 -2533
rect -896 -2635 -862 -2601
rect -815 -2635 -781 -2601
rect -734 -2635 -700 -2601
rect -896 -2703 -862 -2669
rect -815 -2703 -781 -2669
rect -734 -2703 -700 -2669
rect -896 -2771 -862 -2737
rect -815 -2771 -781 -2737
rect -734 -2771 -700 -2737
rect -896 -2839 -862 -2805
rect -815 -2839 -781 -2805
rect -734 -2839 -700 -2805
rect -896 -2907 -862 -2873
rect -815 -2907 -781 -2873
rect -734 -2907 -700 -2873
rect -896 -2975 -862 -2941
rect -815 -2975 -781 -2941
rect -734 -2975 -700 -2941
rect -896 -3043 -862 -3009
rect -815 -3043 -781 -3009
rect -734 -3043 -700 -3009
rect -896 -3111 -862 -3077
rect -815 -3111 -781 -3077
rect -734 -3111 -700 -3077
rect -896 -3179 -862 -3145
rect -815 -3179 -781 -3145
rect -734 -3179 -700 -3145
rect -896 -3247 -862 -3213
rect -815 -3247 -781 -3213
rect -734 -3247 -700 -3213
rect -896 -3315 -862 -3281
rect -815 -3315 -781 -3281
rect -734 -3315 -700 -3281
rect -896 -3383 -862 -3349
rect -815 -3383 -781 -3349
rect -734 -3383 -700 -3349
rect -896 -3451 -862 -3417
rect -815 -3451 -781 -3417
rect -734 -3451 -700 -3417
rect -896 -3519 -862 -3485
rect -815 -3519 -781 -3485
rect -734 -3519 -700 -3485
rect -896 -3587 -862 -3553
rect -815 -3587 -781 -3553
rect -734 -3587 -700 -3553
rect -896 -3655 -862 -3621
rect -815 -3655 -781 -3621
rect -734 -3655 -700 -3621
rect -896 -3723 -862 -3689
rect -815 -3723 -781 -3689
rect -734 -3723 -700 -3689
rect -896 -3791 -862 -3757
rect -815 -3791 -781 -3757
rect -734 -3791 -700 -3757
rect -896 -3859 -862 -3825
rect -815 -3859 -781 -3825
rect -734 -3859 -700 -3825
rect -896 -3927 -862 -3893
rect -815 -3927 -781 -3893
rect -734 -3927 -700 -3893
rect -896 -3995 -862 -3961
rect -815 -3995 -781 -3961
rect -734 -3995 -700 -3961
rect -896 -4063 -862 -4029
rect -815 -4063 -781 -4029
rect -734 -4063 -700 -4029
rect -896 -4131 -862 -4097
rect -815 -4131 -781 -4097
rect -734 -4131 -700 -4097
rect -896 -4199 -862 -4165
rect -815 -4199 -781 -4165
rect -734 -4199 -700 -4165
rect -896 -4267 -862 -4233
rect -815 -4267 -781 -4233
rect -734 -4267 -700 -4233
rect -896 -4335 -862 -4301
rect -815 -4335 -781 -4301
rect -734 -4335 -700 -4301
rect -896 -4403 -862 -4369
rect -815 -4403 -781 -4369
rect -734 -4403 -700 -4369
rect -896 -4471 -862 -4437
rect -815 -4471 -781 -4437
rect -734 -4471 -700 -4437
rect -896 -4539 -862 -4505
rect -815 -4539 -781 -4505
rect -734 -4539 -700 -4505
rect -896 -4607 -862 -4573
rect -815 -4607 -781 -4573
rect -734 -4607 -700 -4573
rect -896 -4675 -862 -4641
rect -815 -4675 -781 -4641
rect -734 -4675 -700 -4641
rect -896 -4743 -862 -4709
rect -815 -4743 -781 -4709
rect -734 -4743 -700 -4709
rect -896 -4811 -862 -4777
rect -815 -4811 -781 -4777
rect -734 -4811 -700 -4777
rect -896 -4879 -862 -4845
rect -815 -4879 -781 -4845
rect -734 -4879 -700 -4845
rect -896 -4947 -862 -4913
rect -815 -4947 -781 -4913
rect -734 -4947 -700 -4913
rect -896 -5015 -862 -4981
rect -815 -5015 -781 -4981
rect -734 -5015 -700 -4981
rect -364 4981 -330 5015
rect -283 4981 -249 5015
rect -202 4981 -168 5015
rect -364 4913 -330 4947
rect -283 4913 -249 4947
rect -202 4913 -168 4947
rect -364 4845 -330 4879
rect -283 4845 -249 4879
rect -202 4845 -168 4879
rect -364 4777 -330 4811
rect -283 4777 -249 4811
rect -202 4777 -168 4811
rect -364 4709 -330 4743
rect -283 4709 -249 4743
rect -202 4709 -168 4743
rect -364 4641 -330 4675
rect -283 4641 -249 4675
rect -202 4641 -168 4675
rect -364 4573 -330 4607
rect -283 4573 -249 4607
rect -202 4573 -168 4607
rect -364 4505 -330 4539
rect -283 4505 -249 4539
rect -202 4505 -168 4539
rect -364 4437 -330 4471
rect -283 4437 -249 4471
rect -202 4437 -168 4471
rect -364 4369 -330 4403
rect -283 4369 -249 4403
rect -202 4369 -168 4403
rect -364 4301 -330 4335
rect -283 4301 -249 4335
rect -202 4301 -168 4335
rect -364 4233 -330 4267
rect -283 4233 -249 4267
rect -202 4233 -168 4267
rect -364 4165 -330 4199
rect -283 4165 -249 4199
rect -202 4165 -168 4199
rect -364 4097 -330 4131
rect -283 4097 -249 4131
rect -202 4097 -168 4131
rect -364 4029 -330 4063
rect -283 4029 -249 4063
rect -202 4029 -168 4063
rect -364 3961 -330 3995
rect -283 3961 -249 3995
rect -202 3961 -168 3995
rect -364 3893 -330 3927
rect -283 3893 -249 3927
rect -202 3893 -168 3927
rect -364 3825 -330 3859
rect -283 3825 -249 3859
rect -202 3825 -168 3859
rect -364 3757 -330 3791
rect -283 3757 -249 3791
rect -202 3757 -168 3791
rect -364 3689 -330 3723
rect -283 3689 -249 3723
rect -202 3689 -168 3723
rect -364 3621 -330 3655
rect -283 3621 -249 3655
rect -202 3621 -168 3655
rect -364 3553 -330 3587
rect -283 3553 -249 3587
rect -202 3553 -168 3587
rect -364 3485 -330 3519
rect -283 3485 -249 3519
rect -202 3485 -168 3519
rect -364 3417 -330 3451
rect -283 3417 -249 3451
rect -202 3417 -168 3451
rect -364 3349 -330 3383
rect -283 3349 -249 3383
rect -202 3349 -168 3383
rect -364 3281 -330 3315
rect -283 3281 -249 3315
rect -202 3281 -168 3315
rect -364 3213 -330 3247
rect -283 3213 -249 3247
rect -202 3213 -168 3247
rect -364 3145 -330 3179
rect -283 3145 -249 3179
rect -202 3145 -168 3179
rect -364 3077 -330 3111
rect -283 3077 -249 3111
rect -202 3077 -168 3111
rect -364 3009 -330 3043
rect -283 3009 -249 3043
rect -202 3009 -168 3043
rect -364 2941 -330 2975
rect -283 2941 -249 2975
rect -202 2941 -168 2975
rect -364 2873 -330 2907
rect -283 2873 -249 2907
rect -202 2873 -168 2907
rect -364 2805 -330 2839
rect -283 2805 -249 2839
rect -202 2805 -168 2839
rect -364 2737 -330 2771
rect -283 2737 -249 2771
rect -202 2737 -168 2771
rect -364 2669 -330 2703
rect -283 2669 -249 2703
rect -202 2669 -168 2703
rect -364 2601 -330 2635
rect -283 2601 -249 2635
rect -202 2601 -168 2635
rect -364 2533 -330 2567
rect -283 2533 -249 2567
rect -202 2533 -168 2567
rect -364 2465 -330 2499
rect -283 2465 -249 2499
rect -202 2465 -168 2499
rect -364 2397 -330 2431
rect -283 2397 -249 2431
rect -202 2397 -168 2431
rect -364 2329 -330 2363
rect -283 2329 -249 2363
rect -202 2329 -168 2363
rect -364 2261 -330 2295
rect -283 2261 -249 2295
rect -202 2261 -168 2295
rect -364 2193 -330 2227
rect -283 2193 -249 2227
rect -202 2193 -168 2227
rect -364 2125 -330 2159
rect -283 2125 -249 2159
rect -202 2125 -168 2159
rect -364 2057 -330 2091
rect -283 2057 -249 2091
rect -202 2057 -168 2091
rect -364 1989 -330 2023
rect -283 1989 -249 2023
rect -202 1989 -168 2023
rect -364 1921 -330 1955
rect -283 1921 -249 1955
rect -202 1921 -168 1955
rect -364 1853 -330 1887
rect -283 1853 -249 1887
rect -202 1853 -168 1887
rect -364 1785 -330 1819
rect -283 1785 -249 1819
rect -202 1785 -168 1819
rect -364 1717 -330 1751
rect -283 1717 -249 1751
rect -202 1717 -168 1751
rect -364 1649 -330 1683
rect -283 1649 -249 1683
rect -202 1649 -168 1683
rect -364 1581 -330 1615
rect -283 1581 -249 1615
rect -202 1581 -168 1615
rect -364 1513 -330 1547
rect -283 1513 -249 1547
rect -202 1513 -168 1547
rect -364 1445 -330 1479
rect -283 1445 -249 1479
rect -202 1445 -168 1479
rect -364 1377 -330 1411
rect -283 1377 -249 1411
rect -202 1377 -168 1411
rect -364 1309 -330 1343
rect -283 1309 -249 1343
rect -202 1309 -168 1343
rect -364 1241 -330 1275
rect -283 1241 -249 1275
rect -202 1241 -168 1275
rect -364 1173 -330 1207
rect -283 1173 -249 1207
rect -202 1173 -168 1207
rect -364 1105 -330 1139
rect -283 1105 -249 1139
rect -202 1105 -168 1139
rect -364 1037 -330 1071
rect -283 1037 -249 1071
rect -202 1037 -168 1071
rect -364 969 -330 1003
rect -283 969 -249 1003
rect -202 969 -168 1003
rect -364 901 -330 935
rect -283 901 -249 935
rect -202 901 -168 935
rect -364 833 -330 867
rect -283 833 -249 867
rect -202 833 -168 867
rect -364 765 -330 799
rect -283 765 -249 799
rect -202 765 -168 799
rect -364 697 -330 731
rect -283 697 -249 731
rect -202 697 -168 731
rect -364 629 -330 663
rect -283 629 -249 663
rect -202 629 -168 663
rect -364 561 -330 595
rect -283 561 -249 595
rect -202 561 -168 595
rect -364 493 -330 527
rect -283 493 -249 527
rect -202 493 -168 527
rect -364 425 -330 459
rect -283 425 -249 459
rect -202 425 -168 459
rect -364 357 -330 391
rect -283 357 -249 391
rect -202 357 -168 391
rect -364 289 -330 323
rect -283 289 -249 323
rect -202 289 -168 323
rect -364 221 -330 255
rect -283 221 -249 255
rect -202 221 -168 255
rect -364 153 -330 187
rect -283 153 -249 187
rect -202 153 -168 187
rect -364 85 -330 119
rect -283 85 -249 119
rect -202 85 -168 119
rect -364 17 -330 51
rect -283 17 -249 51
rect -202 17 -168 51
rect -364 -51 -330 -17
rect -283 -51 -249 -17
rect -202 -51 -168 -17
rect -364 -119 -330 -85
rect -283 -119 -249 -85
rect -202 -119 -168 -85
rect -364 -187 -330 -153
rect -283 -187 -249 -153
rect -202 -187 -168 -153
rect -364 -255 -330 -221
rect -283 -255 -249 -221
rect -202 -255 -168 -221
rect -364 -323 -330 -289
rect -283 -323 -249 -289
rect -202 -323 -168 -289
rect -364 -391 -330 -357
rect -283 -391 -249 -357
rect -202 -391 -168 -357
rect -364 -459 -330 -425
rect -283 -459 -249 -425
rect -202 -459 -168 -425
rect -364 -527 -330 -493
rect -283 -527 -249 -493
rect -202 -527 -168 -493
rect -364 -595 -330 -561
rect -283 -595 -249 -561
rect -202 -595 -168 -561
rect -364 -663 -330 -629
rect -283 -663 -249 -629
rect -202 -663 -168 -629
rect -364 -731 -330 -697
rect -283 -731 -249 -697
rect -202 -731 -168 -697
rect -364 -799 -330 -765
rect -283 -799 -249 -765
rect -202 -799 -168 -765
rect -364 -867 -330 -833
rect -283 -867 -249 -833
rect -202 -867 -168 -833
rect -364 -935 -330 -901
rect -283 -935 -249 -901
rect -202 -935 -168 -901
rect -364 -1003 -330 -969
rect -283 -1003 -249 -969
rect -202 -1003 -168 -969
rect -364 -1071 -330 -1037
rect -283 -1071 -249 -1037
rect -202 -1071 -168 -1037
rect -364 -1139 -330 -1105
rect -283 -1139 -249 -1105
rect -202 -1139 -168 -1105
rect -364 -1207 -330 -1173
rect -283 -1207 -249 -1173
rect -202 -1207 -168 -1173
rect -364 -1275 -330 -1241
rect -283 -1275 -249 -1241
rect -202 -1275 -168 -1241
rect -364 -1343 -330 -1309
rect -283 -1343 -249 -1309
rect -202 -1343 -168 -1309
rect -364 -1411 -330 -1377
rect -283 -1411 -249 -1377
rect -202 -1411 -168 -1377
rect -364 -1479 -330 -1445
rect -283 -1479 -249 -1445
rect -202 -1479 -168 -1445
rect -364 -1547 -330 -1513
rect -283 -1547 -249 -1513
rect -202 -1547 -168 -1513
rect -364 -1615 -330 -1581
rect -283 -1615 -249 -1581
rect -202 -1615 -168 -1581
rect -364 -1683 -330 -1649
rect -283 -1683 -249 -1649
rect -202 -1683 -168 -1649
rect -364 -1751 -330 -1717
rect -283 -1751 -249 -1717
rect -202 -1751 -168 -1717
rect -364 -1819 -330 -1785
rect -283 -1819 -249 -1785
rect -202 -1819 -168 -1785
rect -364 -1887 -330 -1853
rect -283 -1887 -249 -1853
rect -202 -1887 -168 -1853
rect -364 -1955 -330 -1921
rect -283 -1955 -249 -1921
rect -202 -1955 -168 -1921
rect -364 -2023 -330 -1989
rect -283 -2023 -249 -1989
rect -202 -2023 -168 -1989
rect -364 -2091 -330 -2057
rect -283 -2091 -249 -2057
rect -202 -2091 -168 -2057
rect -364 -2159 -330 -2125
rect -283 -2159 -249 -2125
rect -202 -2159 -168 -2125
rect -364 -2227 -330 -2193
rect -283 -2227 -249 -2193
rect -202 -2227 -168 -2193
rect -364 -2295 -330 -2261
rect -283 -2295 -249 -2261
rect -202 -2295 -168 -2261
rect -364 -2363 -330 -2329
rect -283 -2363 -249 -2329
rect -202 -2363 -168 -2329
rect -364 -2431 -330 -2397
rect -283 -2431 -249 -2397
rect -202 -2431 -168 -2397
rect -364 -2499 -330 -2465
rect -283 -2499 -249 -2465
rect -202 -2499 -168 -2465
rect -364 -2567 -330 -2533
rect -283 -2567 -249 -2533
rect -202 -2567 -168 -2533
rect -364 -2635 -330 -2601
rect -283 -2635 -249 -2601
rect -202 -2635 -168 -2601
rect -364 -2703 -330 -2669
rect -283 -2703 -249 -2669
rect -202 -2703 -168 -2669
rect -364 -2771 -330 -2737
rect -283 -2771 -249 -2737
rect -202 -2771 -168 -2737
rect -364 -2839 -330 -2805
rect -283 -2839 -249 -2805
rect -202 -2839 -168 -2805
rect -364 -2907 -330 -2873
rect -283 -2907 -249 -2873
rect -202 -2907 -168 -2873
rect -364 -2975 -330 -2941
rect -283 -2975 -249 -2941
rect -202 -2975 -168 -2941
rect -364 -3043 -330 -3009
rect -283 -3043 -249 -3009
rect -202 -3043 -168 -3009
rect -364 -3111 -330 -3077
rect -283 -3111 -249 -3077
rect -202 -3111 -168 -3077
rect -364 -3179 -330 -3145
rect -283 -3179 -249 -3145
rect -202 -3179 -168 -3145
rect -364 -3247 -330 -3213
rect -283 -3247 -249 -3213
rect -202 -3247 -168 -3213
rect -364 -3315 -330 -3281
rect -283 -3315 -249 -3281
rect -202 -3315 -168 -3281
rect -364 -3383 -330 -3349
rect -283 -3383 -249 -3349
rect -202 -3383 -168 -3349
rect -364 -3451 -330 -3417
rect -283 -3451 -249 -3417
rect -202 -3451 -168 -3417
rect -364 -3519 -330 -3485
rect -283 -3519 -249 -3485
rect -202 -3519 -168 -3485
rect -364 -3587 -330 -3553
rect -283 -3587 -249 -3553
rect -202 -3587 -168 -3553
rect -364 -3655 -330 -3621
rect -283 -3655 -249 -3621
rect -202 -3655 -168 -3621
rect -364 -3723 -330 -3689
rect -283 -3723 -249 -3689
rect -202 -3723 -168 -3689
rect -364 -3791 -330 -3757
rect -283 -3791 -249 -3757
rect -202 -3791 -168 -3757
rect -364 -3859 -330 -3825
rect -283 -3859 -249 -3825
rect -202 -3859 -168 -3825
rect -364 -3927 -330 -3893
rect -283 -3927 -249 -3893
rect -202 -3927 -168 -3893
rect -364 -3995 -330 -3961
rect -283 -3995 -249 -3961
rect -202 -3995 -168 -3961
rect -364 -4063 -330 -4029
rect -283 -4063 -249 -4029
rect -202 -4063 -168 -4029
rect -364 -4131 -330 -4097
rect -283 -4131 -249 -4097
rect -202 -4131 -168 -4097
rect -364 -4199 -330 -4165
rect -283 -4199 -249 -4165
rect -202 -4199 -168 -4165
rect -364 -4267 -330 -4233
rect -283 -4267 -249 -4233
rect -202 -4267 -168 -4233
rect -364 -4335 -330 -4301
rect -283 -4335 -249 -4301
rect -202 -4335 -168 -4301
rect -364 -4403 -330 -4369
rect -283 -4403 -249 -4369
rect -202 -4403 -168 -4369
rect -364 -4471 -330 -4437
rect -283 -4471 -249 -4437
rect -202 -4471 -168 -4437
rect -364 -4539 -330 -4505
rect -283 -4539 -249 -4505
rect -202 -4539 -168 -4505
rect -364 -4607 -330 -4573
rect -283 -4607 -249 -4573
rect -202 -4607 -168 -4573
rect -364 -4675 -330 -4641
rect -283 -4675 -249 -4641
rect -202 -4675 -168 -4641
rect -364 -4743 -330 -4709
rect -283 -4743 -249 -4709
rect -202 -4743 -168 -4709
rect -364 -4811 -330 -4777
rect -283 -4811 -249 -4777
rect -202 -4811 -168 -4777
rect -364 -4879 -330 -4845
rect -283 -4879 -249 -4845
rect -202 -4879 -168 -4845
rect -364 -4947 -330 -4913
rect -283 -4947 -249 -4913
rect -202 -4947 -168 -4913
rect -364 -5015 -330 -4981
rect -283 -5015 -249 -4981
rect -202 -5015 -168 -4981
rect 168 4981 202 5015
rect 249 4981 283 5015
rect 330 4981 364 5015
rect 168 4913 202 4947
rect 249 4913 283 4947
rect 330 4913 364 4947
rect 168 4845 202 4879
rect 249 4845 283 4879
rect 330 4845 364 4879
rect 168 4777 202 4811
rect 249 4777 283 4811
rect 330 4777 364 4811
rect 168 4709 202 4743
rect 249 4709 283 4743
rect 330 4709 364 4743
rect 168 4641 202 4675
rect 249 4641 283 4675
rect 330 4641 364 4675
rect 168 4573 202 4607
rect 249 4573 283 4607
rect 330 4573 364 4607
rect 168 4505 202 4539
rect 249 4505 283 4539
rect 330 4505 364 4539
rect 168 4437 202 4471
rect 249 4437 283 4471
rect 330 4437 364 4471
rect 168 4369 202 4403
rect 249 4369 283 4403
rect 330 4369 364 4403
rect 168 4301 202 4335
rect 249 4301 283 4335
rect 330 4301 364 4335
rect 168 4233 202 4267
rect 249 4233 283 4267
rect 330 4233 364 4267
rect 168 4165 202 4199
rect 249 4165 283 4199
rect 330 4165 364 4199
rect 168 4097 202 4131
rect 249 4097 283 4131
rect 330 4097 364 4131
rect 168 4029 202 4063
rect 249 4029 283 4063
rect 330 4029 364 4063
rect 168 3961 202 3995
rect 249 3961 283 3995
rect 330 3961 364 3995
rect 168 3893 202 3927
rect 249 3893 283 3927
rect 330 3893 364 3927
rect 168 3825 202 3859
rect 249 3825 283 3859
rect 330 3825 364 3859
rect 168 3757 202 3791
rect 249 3757 283 3791
rect 330 3757 364 3791
rect 168 3689 202 3723
rect 249 3689 283 3723
rect 330 3689 364 3723
rect 168 3621 202 3655
rect 249 3621 283 3655
rect 330 3621 364 3655
rect 168 3553 202 3587
rect 249 3553 283 3587
rect 330 3553 364 3587
rect 168 3485 202 3519
rect 249 3485 283 3519
rect 330 3485 364 3519
rect 168 3417 202 3451
rect 249 3417 283 3451
rect 330 3417 364 3451
rect 168 3349 202 3383
rect 249 3349 283 3383
rect 330 3349 364 3383
rect 168 3281 202 3315
rect 249 3281 283 3315
rect 330 3281 364 3315
rect 168 3213 202 3247
rect 249 3213 283 3247
rect 330 3213 364 3247
rect 168 3145 202 3179
rect 249 3145 283 3179
rect 330 3145 364 3179
rect 168 3077 202 3111
rect 249 3077 283 3111
rect 330 3077 364 3111
rect 168 3009 202 3043
rect 249 3009 283 3043
rect 330 3009 364 3043
rect 168 2941 202 2975
rect 249 2941 283 2975
rect 330 2941 364 2975
rect 168 2873 202 2907
rect 249 2873 283 2907
rect 330 2873 364 2907
rect 168 2805 202 2839
rect 249 2805 283 2839
rect 330 2805 364 2839
rect 168 2737 202 2771
rect 249 2737 283 2771
rect 330 2737 364 2771
rect 168 2669 202 2703
rect 249 2669 283 2703
rect 330 2669 364 2703
rect 168 2601 202 2635
rect 249 2601 283 2635
rect 330 2601 364 2635
rect 168 2533 202 2567
rect 249 2533 283 2567
rect 330 2533 364 2567
rect 168 2465 202 2499
rect 249 2465 283 2499
rect 330 2465 364 2499
rect 168 2397 202 2431
rect 249 2397 283 2431
rect 330 2397 364 2431
rect 168 2329 202 2363
rect 249 2329 283 2363
rect 330 2329 364 2363
rect 168 2261 202 2295
rect 249 2261 283 2295
rect 330 2261 364 2295
rect 168 2193 202 2227
rect 249 2193 283 2227
rect 330 2193 364 2227
rect 168 2125 202 2159
rect 249 2125 283 2159
rect 330 2125 364 2159
rect 168 2057 202 2091
rect 249 2057 283 2091
rect 330 2057 364 2091
rect 168 1989 202 2023
rect 249 1989 283 2023
rect 330 1989 364 2023
rect 168 1921 202 1955
rect 249 1921 283 1955
rect 330 1921 364 1955
rect 168 1853 202 1887
rect 249 1853 283 1887
rect 330 1853 364 1887
rect 168 1785 202 1819
rect 249 1785 283 1819
rect 330 1785 364 1819
rect 168 1717 202 1751
rect 249 1717 283 1751
rect 330 1717 364 1751
rect 168 1649 202 1683
rect 249 1649 283 1683
rect 330 1649 364 1683
rect 168 1581 202 1615
rect 249 1581 283 1615
rect 330 1581 364 1615
rect 168 1513 202 1547
rect 249 1513 283 1547
rect 330 1513 364 1547
rect 168 1445 202 1479
rect 249 1445 283 1479
rect 330 1445 364 1479
rect 168 1377 202 1411
rect 249 1377 283 1411
rect 330 1377 364 1411
rect 168 1309 202 1343
rect 249 1309 283 1343
rect 330 1309 364 1343
rect 168 1241 202 1275
rect 249 1241 283 1275
rect 330 1241 364 1275
rect 168 1173 202 1207
rect 249 1173 283 1207
rect 330 1173 364 1207
rect 168 1105 202 1139
rect 249 1105 283 1139
rect 330 1105 364 1139
rect 168 1037 202 1071
rect 249 1037 283 1071
rect 330 1037 364 1071
rect 168 969 202 1003
rect 249 969 283 1003
rect 330 969 364 1003
rect 168 901 202 935
rect 249 901 283 935
rect 330 901 364 935
rect 168 833 202 867
rect 249 833 283 867
rect 330 833 364 867
rect 168 765 202 799
rect 249 765 283 799
rect 330 765 364 799
rect 168 697 202 731
rect 249 697 283 731
rect 330 697 364 731
rect 168 629 202 663
rect 249 629 283 663
rect 330 629 364 663
rect 168 561 202 595
rect 249 561 283 595
rect 330 561 364 595
rect 168 493 202 527
rect 249 493 283 527
rect 330 493 364 527
rect 168 425 202 459
rect 249 425 283 459
rect 330 425 364 459
rect 168 357 202 391
rect 249 357 283 391
rect 330 357 364 391
rect 168 289 202 323
rect 249 289 283 323
rect 330 289 364 323
rect 168 221 202 255
rect 249 221 283 255
rect 330 221 364 255
rect 168 153 202 187
rect 249 153 283 187
rect 330 153 364 187
rect 168 85 202 119
rect 249 85 283 119
rect 330 85 364 119
rect 168 17 202 51
rect 249 17 283 51
rect 330 17 364 51
rect 168 -51 202 -17
rect 249 -51 283 -17
rect 330 -51 364 -17
rect 168 -119 202 -85
rect 249 -119 283 -85
rect 330 -119 364 -85
rect 168 -187 202 -153
rect 249 -187 283 -153
rect 330 -187 364 -153
rect 168 -255 202 -221
rect 249 -255 283 -221
rect 330 -255 364 -221
rect 168 -323 202 -289
rect 249 -323 283 -289
rect 330 -323 364 -289
rect 168 -391 202 -357
rect 249 -391 283 -357
rect 330 -391 364 -357
rect 168 -459 202 -425
rect 249 -459 283 -425
rect 330 -459 364 -425
rect 168 -527 202 -493
rect 249 -527 283 -493
rect 330 -527 364 -493
rect 168 -595 202 -561
rect 249 -595 283 -561
rect 330 -595 364 -561
rect 168 -663 202 -629
rect 249 -663 283 -629
rect 330 -663 364 -629
rect 168 -731 202 -697
rect 249 -731 283 -697
rect 330 -731 364 -697
rect 168 -799 202 -765
rect 249 -799 283 -765
rect 330 -799 364 -765
rect 168 -867 202 -833
rect 249 -867 283 -833
rect 330 -867 364 -833
rect 168 -935 202 -901
rect 249 -935 283 -901
rect 330 -935 364 -901
rect 168 -1003 202 -969
rect 249 -1003 283 -969
rect 330 -1003 364 -969
rect 168 -1071 202 -1037
rect 249 -1071 283 -1037
rect 330 -1071 364 -1037
rect 168 -1139 202 -1105
rect 249 -1139 283 -1105
rect 330 -1139 364 -1105
rect 168 -1207 202 -1173
rect 249 -1207 283 -1173
rect 330 -1207 364 -1173
rect 168 -1275 202 -1241
rect 249 -1275 283 -1241
rect 330 -1275 364 -1241
rect 168 -1343 202 -1309
rect 249 -1343 283 -1309
rect 330 -1343 364 -1309
rect 168 -1411 202 -1377
rect 249 -1411 283 -1377
rect 330 -1411 364 -1377
rect 168 -1479 202 -1445
rect 249 -1479 283 -1445
rect 330 -1479 364 -1445
rect 168 -1547 202 -1513
rect 249 -1547 283 -1513
rect 330 -1547 364 -1513
rect 168 -1615 202 -1581
rect 249 -1615 283 -1581
rect 330 -1615 364 -1581
rect 168 -1683 202 -1649
rect 249 -1683 283 -1649
rect 330 -1683 364 -1649
rect 168 -1751 202 -1717
rect 249 -1751 283 -1717
rect 330 -1751 364 -1717
rect 168 -1819 202 -1785
rect 249 -1819 283 -1785
rect 330 -1819 364 -1785
rect 168 -1887 202 -1853
rect 249 -1887 283 -1853
rect 330 -1887 364 -1853
rect 168 -1955 202 -1921
rect 249 -1955 283 -1921
rect 330 -1955 364 -1921
rect 168 -2023 202 -1989
rect 249 -2023 283 -1989
rect 330 -2023 364 -1989
rect 168 -2091 202 -2057
rect 249 -2091 283 -2057
rect 330 -2091 364 -2057
rect 168 -2159 202 -2125
rect 249 -2159 283 -2125
rect 330 -2159 364 -2125
rect 168 -2227 202 -2193
rect 249 -2227 283 -2193
rect 330 -2227 364 -2193
rect 168 -2295 202 -2261
rect 249 -2295 283 -2261
rect 330 -2295 364 -2261
rect 168 -2363 202 -2329
rect 249 -2363 283 -2329
rect 330 -2363 364 -2329
rect 168 -2431 202 -2397
rect 249 -2431 283 -2397
rect 330 -2431 364 -2397
rect 168 -2499 202 -2465
rect 249 -2499 283 -2465
rect 330 -2499 364 -2465
rect 168 -2567 202 -2533
rect 249 -2567 283 -2533
rect 330 -2567 364 -2533
rect 168 -2635 202 -2601
rect 249 -2635 283 -2601
rect 330 -2635 364 -2601
rect 168 -2703 202 -2669
rect 249 -2703 283 -2669
rect 330 -2703 364 -2669
rect 168 -2771 202 -2737
rect 249 -2771 283 -2737
rect 330 -2771 364 -2737
rect 168 -2839 202 -2805
rect 249 -2839 283 -2805
rect 330 -2839 364 -2805
rect 168 -2907 202 -2873
rect 249 -2907 283 -2873
rect 330 -2907 364 -2873
rect 168 -2975 202 -2941
rect 249 -2975 283 -2941
rect 330 -2975 364 -2941
rect 168 -3043 202 -3009
rect 249 -3043 283 -3009
rect 330 -3043 364 -3009
rect 168 -3111 202 -3077
rect 249 -3111 283 -3077
rect 330 -3111 364 -3077
rect 168 -3179 202 -3145
rect 249 -3179 283 -3145
rect 330 -3179 364 -3145
rect 168 -3247 202 -3213
rect 249 -3247 283 -3213
rect 330 -3247 364 -3213
rect 168 -3315 202 -3281
rect 249 -3315 283 -3281
rect 330 -3315 364 -3281
rect 168 -3383 202 -3349
rect 249 -3383 283 -3349
rect 330 -3383 364 -3349
rect 168 -3451 202 -3417
rect 249 -3451 283 -3417
rect 330 -3451 364 -3417
rect 168 -3519 202 -3485
rect 249 -3519 283 -3485
rect 330 -3519 364 -3485
rect 168 -3587 202 -3553
rect 249 -3587 283 -3553
rect 330 -3587 364 -3553
rect 168 -3655 202 -3621
rect 249 -3655 283 -3621
rect 330 -3655 364 -3621
rect 168 -3723 202 -3689
rect 249 -3723 283 -3689
rect 330 -3723 364 -3689
rect 168 -3791 202 -3757
rect 249 -3791 283 -3757
rect 330 -3791 364 -3757
rect 168 -3859 202 -3825
rect 249 -3859 283 -3825
rect 330 -3859 364 -3825
rect 168 -3927 202 -3893
rect 249 -3927 283 -3893
rect 330 -3927 364 -3893
rect 168 -3995 202 -3961
rect 249 -3995 283 -3961
rect 330 -3995 364 -3961
rect 168 -4063 202 -4029
rect 249 -4063 283 -4029
rect 330 -4063 364 -4029
rect 168 -4131 202 -4097
rect 249 -4131 283 -4097
rect 330 -4131 364 -4097
rect 168 -4199 202 -4165
rect 249 -4199 283 -4165
rect 330 -4199 364 -4165
rect 168 -4267 202 -4233
rect 249 -4267 283 -4233
rect 330 -4267 364 -4233
rect 168 -4335 202 -4301
rect 249 -4335 283 -4301
rect 330 -4335 364 -4301
rect 168 -4403 202 -4369
rect 249 -4403 283 -4369
rect 330 -4403 364 -4369
rect 168 -4471 202 -4437
rect 249 -4471 283 -4437
rect 330 -4471 364 -4437
rect 168 -4539 202 -4505
rect 249 -4539 283 -4505
rect 330 -4539 364 -4505
rect 168 -4607 202 -4573
rect 249 -4607 283 -4573
rect 330 -4607 364 -4573
rect 168 -4675 202 -4641
rect 249 -4675 283 -4641
rect 330 -4675 364 -4641
rect 168 -4743 202 -4709
rect 249 -4743 283 -4709
rect 330 -4743 364 -4709
rect 168 -4811 202 -4777
rect 249 -4811 283 -4777
rect 330 -4811 364 -4777
rect 168 -4879 202 -4845
rect 249 -4879 283 -4845
rect 330 -4879 364 -4845
rect 168 -4947 202 -4913
rect 249 -4947 283 -4913
rect 330 -4947 364 -4913
rect 168 -5015 202 -4981
rect 249 -5015 283 -4981
rect 330 -5015 364 -4981
rect 700 4981 734 5015
rect 781 4981 815 5015
rect 862 4981 896 5015
rect 700 4913 734 4947
rect 781 4913 815 4947
rect 862 4913 896 4947
rect 700 4845 734 4879
rect 781 4845 815 4879
rect 862 4845 896 4879
rect 700 4777 734 4811
rect 781 4777 815 4811
rect 862 4777 896 4811
rect 700 4709 734 4743
rect 781 4709 815 4743
rect 862 4709 896 4743
rect 700 4641 734 4675
rect 781 4641 815 4675
rect 862 4641 896 4675
rect 700 4573 734 4607
rect 781 4573 815 4607
rect 862 4573 896 4607
rect 700 4505 734 4539
rect 781 4505 815 4539
rect 862 4505 896 4539
rect 700 4437 734 4471
rect 781 4437 815 4471
rect 862 4437 896 4471
rect 700 4369 734 4403
rect 781 4369 815 4403
rect 862 4369 896 4403
rect 700 4301 734 4335
rect 781 4301 815 4335
rect 862 4301 896 4335
rect 700 4233 734 4267
rect 781 4233 815 4267
rect 862 4233 896 4267
rect 700 4165 734 4199
rect 781 4165 815 4199
rect 862 4165 896 4199
rect 700 4097 734 4131
rect 781 4097 815 4131
rect 862 4097 896 4131
rect 700 4029 734 4063
rect 781 4029 815 4063
rect 862 4029 896 4063
rect 700 3961 734 3995
rect 781 3961 815 3995
rect 862 3961 896 3995
rect 700 3893 734 3927
rect 781 3893 815 3927
rect 862 3893 896 3927
rect 700 3825 734 3859
rect 781 3825 815 3859
rect 862 3825 896 3859
rect 700 3757 734 3791
rect 781 3757 815 3791
rect 862 3757 896 3791
rect 700 3689 734 3723
rect 781 3689 815 3723
rect 862 3689 896 3723
rect 700 3621 734 3655
rect 781 3621 815 3655
rect 862 3621 896 3655
rect 700 3553 734 3587
rect 781 3553 815 3587
rect 862 3553 896 3587
rect 700 3485 734 3519
rect 781 3485 815 3519
rect 862 3485 896 3519
rect 700 3417 734 3451
rect 781 3417 815 3451
rect 862 3417 896 3451
rect 700 3349 734 3383
rect 781 3349 815 3383
rect 862 3349 896 3383
rect 700 3281 734 3315
rect 781 3281 815 3315
rect 862 3281 896 3315
rect 700 3213 734 3247
rect 781 3213 815 3247
rect 862 3213 896 3247
rect 700 3145 734 3179
rect 781 3145 815 3179
rect 862 3145 896 3179
rect 700 3077 734 3111
rect 781 3077 815 3111
rect 862 3077 896 3111
rect 700 3009 734 3043
rect 781 3009 815 3043
rect 862 3009 896 3043
rect 700 2941 734 2975
rect 781 2941 815 2975
rect 862 2941 896 2975
rect 700 2873 734 2907
rect 781 2873 815 2907
rect 862 2873 896 2907
rect 700 2805 734 2839
rect 781 2805 815 2839
rect 862 2805 896 2839
rect 700 2737 734 2771
rect 781 2737 815 2771
rect 862 2737 896 2771
rect 700 2669 734 2703
rect 781 2669 815 2703
rect 862 2669 896 2703
rect 700 2601 734 2635
rect 781 2601 815 2635
rect 862 2601 896 2635
rect 700 2533 734 2567
rect 781 2533 815 2567
rect 862 2533 896 2567
rect 700 2465 734 2499
rect 781 2465 815 2499
rect 862 2465 896 2499
rect 700 2397 734 2431
rect 781 2397 815 2431
rect 862 2397 896 2431
rect 700 2329 734 2363
rect 781 2329 815 2363
rect 862 2329 896 2363
rect 700 2261 734 2295
rect 781 2261 815 2295
rect 862 2261 896 2295
rect 700 2193 734 2227
rect 781 2193 815 2227
rect 862 2193 896 2227
rect 700 2125 734 2159
rect 781 2125 815 2159
rect 862 2125 896 2159
rect 700 2057 734 2091
rect 781 2057 815 2091
rect 862 2057 896 2091
rect 700 1989 734 2023
rect 781 1989 815 2023
rect 862 1989 896 2023
rect 700 1921 734 1955
rect 781 1921 815 1955
rect 862 1921 896 1955
rect 700 1853 734 1887
rect 781 1853 815 1887
rect 862 1853 896 1887
rect 700 1785 734 1819
rect 781 1785 815 1819
rect 862 1785 896 1819
rect 700 1717 734 1751
rect 781 1717 815 1751
rect 862 1717 896 1751
rect 700 1649 734 1683
rect 781 1649 815 1683
rect 862 1649 896 1683
rect 700 1581 734 1615
rect 781 1581 815 1615
rect 862 1581 896 1615
rect 700 1513 734 1547
rect 781 1513 815 1547
rect 862 1513 896 1547
rect 700 1445 734 1479
rect 781 1445 815 1479
rect 862 1445 896 1479
rect 700 1377 734 1411
rect 781 1377 815 1411
rect 862 1377 896 1411
rect 700 1309 734 1343
rect 781 1309 815 1343
rect 862 1309 896 1343
rect 700 1241 734 1275
rect 781 1241 815 1275
rect 862 1241 896 1275
rect 700 1173 734 1207
rect 781 1173 815 1207
rect 862 1173 896 1207
rect 700 1105 734 1139
rect 781 1105 815 1139
rect 862 1105 896 1139
rect 700 1037 734 1071
rect 781 1037 815 1071
rect 862 1037 896 1071
rect 700 969 734 1003
rect 781 969 815 1003
rect 862 969 896 1003
rect 700 901 734 935
rect 781 901 815 935
rect 862 901 896 935
rect 700 833 734 867
rect 781 833 815 867
rect 862 833 896 867
rect 700 765 734 799
rect 781 765 815 799
rect 862 765 896 799
rect 700 697 734 731
rect 781 697 815 731
rect 862 697 896 731
rect 700 629 734 663
rect 781 629 815 663
rect 862 629 896 663
rect 700 561 734 595
rect 781 561 815 595
rect 862 561 896 595
rect 700 493 734 527
rect 781 493 815 527
rect 862 493 896 527
rect 700 425 734 459
rect 781 425 815 459
rect 862 425 896 459
rect 700 357 734 391
rect 781 357 815 391
rect 862 357 896 391
rect 700 289 734 323
rect 781 289 815 323
rect 862 289 896 323
rect 700 221 734 255
rect 781 221 815 255
rect 862 221 896 255
rect 700 153 734 187
rect 781 153 815 187
rect 862 153 896 187
rect 700 85 734 119
rect 781 85 815 119
rect 862 85 896 119
rect 700 17 734 51
rect 781 17 815 51
rect 862 17 896 51
rect 700 -51 734 -17
rect 781 -51 815 -17
rect 862 -51 896 -17
rect 700 -119 734 -85
rect 781 -119 815 -85
rect 862 -119 896 -85
rect 700 -187 734 -153
rect 781 -187 815 -153
rect 862 -187 896 -153
rect 700 -255 734 -221
rect 781 -255 815 -221
rect 862 -255 896 -221
rect 700 -323 734 -289
rect 781 -323 815 -289
rect 862 -323 896 -289
rect 700 -391 734 -357
rect 781 -391 815 -357
rect 862 -391 896 -357
rect 700 -459 734 -425
rect 781 -459 815 -425
rect 862 -459 896 -425
rect 700 -527 734 -493
rect 781 -527 815 -493
rect 862 -527 896 -493
rect 700 -595 734 -561
rect 781 -595 815 -561
rect 862 -595 896 -561
rect 700 -663 734 -629
rect 781 -663 815 -629
rect 862 -663 896 -629
rect 700 -731 734 -697
rect 781 -731 815 -697
rect 862 -731 896 -697
rect 700 -799 734 -765
rect 781 -799 815 -765
rect 862 -799 896 -765
rect 700 -867 734 -833
rect 781 -867 815 -833
rect 862 -867 896 -833
rect 700 -935 734 -901
rect 781 -935 815 -901
rect 862 -935 896 -901
rect 700 -1003 734 -969
rect 781 -1003 815 -969
rect 862 -1003 896 -969
rect 700 -1071 734 -1037
rect 781 -1071 815 -1037
rect 862 -1071 896 -1037
rect 700 -1139 734 -1105
rect 781 -1139 815 -1105
rect 862 -1139 896 -1105
rect 700 -1207 734 -1173
rect 781 -1207 815 -1173
rect 862 -1207 896 -1173
rect 700 -1275 734 -1241
rect 781 -1275 815 -1241
rect 862 -1275 896 -1241
rect 700 -1343 734 -1309
rect 781 -1343 815 -1309
rect 862 -1343 896 -1309
rect 700 -1411 734 -1377
rect 781 -1411 815 -1377
rect 862 -1411 896 -1377
rect 700 -1479 734 -1445
rect 781 -1479 815 -1445
rect 862 -1479 896 -1445
rect 700 -1547 734 -1513
rect 781 -1547 815 -1513
rect 862 -1547 896 -1513
rect 700 -1615 734 -1581
rect 781 -1615 815 -1581
rect 862 -1615 896 -1581
rect 700 -1683 734 -1649
rect 781 -1683 815 -1649
rect 862 -1683 896 -1649
rect 700 -1751 734 -1717
rect 781 -1751 815 -1717
rect 862 -1751 896 -1717
rect 700 -1819 734 -1785
rect 781 -1819 815 -1785
rect 862 -1819 896 -1785
rect 700 -1887 734 -1853
rect 781 -1887 815 -1853
rect 862 -1887 896 -1853
rect 700 -1955 734 -1921
rect 781 -1955 815 -1921
rect 862 -1955 896 -1921
rect 700 -2023 734 -1989
rect 781 -2023 815 -1989
rect 862 -2023 896 -1989
rect 700 -2091 734 -2057
rect 781 -2091 815 -2057
rect 862 -2091 896 -2057
rect 700 -2159 734 -2125
rect 781 -2159 815 -2125
rect 862 -2159 896 -2125
rect 700 -2227 734 -2193
rect 781 -2227 815 -2193
rect 862 -2227 896 -2193
rect 700 -2295 734 -2261
rect 781 -2295 815 -2261
rect 862 -2295 896 -2261
rect 700 -2363 734 -2329
rect 781 -2363 815 -2329
rect 862 -2363 896 -2329
rect 700 -2431 734 -2397
rect 781 -2431 815 -2397
rect 862 -2431 896 -2397
rect 700 -2499 734 -2465
rect 781 -2499 815 -2465
rect 862 -2499 896 -2465
rect 700 -2567 734 -2533
rect 781 -2567 815 -2533
rect 862 -2567 896 -2533
rect 700 -2635 734 -2601
rect 781 -2635 815 -2601
rect 862 -2635 896 -2601
rect 700 -2703 734 -2669
rect 781 -2703 815 -2669
rect 862 -2703 896 -2669
rect 700 -2771 734 -2737
rect 781 -2771 815 -2737
rect 862 -2771 896 -2737
rect 700 -2839 734 -2805
rect 781 -2839 815 -2805
rect 862 -2839 896 -2805
rect 700 -2907 734 -2873
rect 781 -2907 815 -2873
rect 862 -2907 896 -2873
rect 700 -2975 734 -2941
rect 781 -2975 815 -2941
rect 862 -2975 896 -2941
rect 700 -3043 734 -3009
rect 781 -3043 815 -3009
rect 862 -3043 896 -3009
rect 700 -3111 734 -3077
rect 781 -3111 815 -3077
rect 862 -3111 896 -3077
rect 700 -3179 734 -3145
rect 781 -3179 815 -3145
rect 862 -3179 896 -3145
rect 700 -3247 734 -3213
rect 781 -3247 815 -3213
rect 862 -3247 896 -3213
rect 700 -3315 734 -3281
rect 781 -3315 815 -3281
rect 862 -3315 896 -3281
rect 700 -3383 734 -3349
rect 781 -3383 815 -3349
rect 862 -3383 896 -3349
rect 700 -3451 734 -3417
rect 781 -3451 815 -3417
rect 862 -3451 896 -3417
rect 700 -3519 734 -3485
rect 781 -3519 815 -3485
rect 862 -3519 896 -3485
rect 700 -3587 734 -3553
rect 781 -3587 815 -3553
rect 862 -3587 896 -3553
rect 700 -3655 734 -3621
rect 781 -3655 815 -3621
rect 862 -3655 896 -3621
rect 700 -3723 734 -3689
rect 781 -3723 815 -3689
rect 862 -3723 896 -3689
rect 700 -3791 734 -3757
rect 781 -3791 815 -3757
rect 862 -3791 896 -3757
rect 700 -3859 734 -3825
rect 781 -3859 815 -3825
rect 862 -3859 896 -3825
rect 700 -3927 734 -3893
rect 781 -3927 815 -3893
rect 862 -3927 896 -3893
rect 700 -3995 734 -3961
rect 781 -3995 815 -3961
rect 862 -3995 896 -3961
rect 700 -4063 734 -4029
rect 781 -4063 815 -4029
rect 862 -4063 896 -4029
rect 700 -4131 734 -4097
rect 781 -4131 815 -4097
rect 862 -4131 896 -4097
rect 700 -4199 734 -4165
rect 781 -4199 815 -4165
rect 862 -4199 896 -4165
rect 700 -4267 734 -4233
rect 781 -4267 815 -4233
rect 862 -4267 896 -4233
rect 700 -4335 734 -4301
rect 781 -4335 815 -4301
rect 862 -4335 896 -4301
rect 700 -4403 734 -4369
rect 781 -4403 815 -4369
rect 862 -4403 896 -4369
rect 700 -4471 734 -4437
rect 781 -4471 815 -4437
rect 862 -4471 896 -4437
rect 700 -4539 734 -4505
rect 781 -4539 815 -4505
rect 862 -4539 896 -4505
rect 700 -4607 734 -4573
rect 781 -4607 815 -4573
rect 862 -4607 896 -4573
rect 700 -4675 734 -4641
rect 781 -4675 815 -4641
rect 862 -4675 896 -4641
rect 700 -4743 734 -4709
rect 781 -4743 815 -4709
rect 862 -4743 896 -4709
rect 700 -4811 734 -4777
rect 781 -4811 815 -4777
rect 862 -4811 896 -4777
rect 700 -4879 734 -4845
rect 781 -4879 815 -4845
rect 862 -4879 896 -4845
rect 700 -4947 734 -4913
rect 781 -4947 815 -4913
rect 862 -4947 896 -4913
rect 700 -5015 734 -4981
rect 781 -5015 815 -4981
rect 862 -5015 896 -4981
rect 1232 4981 1266 5015
rect 1232 4913 1266 4947
rect 1232 4845 1266 4879
rect 1232 4777 1266 4811
rect 1232 4709 1266 4743
rect 1232 4641 1266 4675
rect 1232 4573 1266 4607
rect 1232 4505 1266 4539
rect 1232 4437 1266 4471
rect 1232 4369 1266 4403
rect 1232 4301 1266 4335
rect 1232 4233 1266 4267
rect 1232 4165 1266 4199
rect 1232 4097 1266 4131
rect 1232 4029 1266 4063
rect 1232 3961 1266 3995
rect 1232 3893 1266 3927
rect 1232 3825 1266 3859
rect 1232 3757 1266 3791
rect 1232 3689 1266 3723
rect 1232 3621 1266 3655
rect 1232 3553 1266 3587
rect 1232 3485 1266 3519
rect 1232 3417 1266 3451
rect 1232 3349 1266 3383
rect 1232 3281 1266 3315
rect 1232 3213 1266 3247
rect 1232 3145 1266 3179
rect 1232 3077 1266 3111
rect 1232 3009 1266 3043
rect 1232 2941 1266 2975
rect 1232 2873 1266 2907
rect 1232 2805 1266 2839
rect 1232 2737 1266 2771
rect 1232 2669 1266 2703
rect 1232 2601 1266 2635
rect 1232 2533 1266 2567
rect 1232 2465 1266 2499
rect 1232 2397 1266 2431
rect 1232 2329 1266 2363
rect 1232 2261 1266 2295
rect 1232 2193 1266 2227
rect 1232 2125 1266 2159
rect 1232 2057 1266 2091
rect 1232 1989 1266 2023
rect 1232 1921 1266 1955
rect 1232 1853 1266 1887
rect 1232 1785 1266 1819
rect 1232 1717 1266 1751
rect 1232 1649 1266 1683
rect 1232 1581 1266 1615
rect 1232 1513 1266 1547
rect 1232 1445 1266 1479
rect 1232 1377 1266 1411
rect 1232 1309 1266 1343
rect 1232 1241 1266 1275
rect 1232 1173 1266 1207
rect 1232 1105 1266 1139
rect 1232 1037 1266 1071
rect 1232 969 1266 1003
rect 1232 901 1266 935
rect 1232 833 1266 867
rect 1232 765 1266 799
rect 1232 697 1266 731
rect 1232 629 1266 663
rect 1232 561 1266 595
rect 1232 493 1266 527
rect 1232 425 1266 459
rect 1232 357 1266 391
rect 1232 289 1266 323
rect 1232 221 1266 255
rect 1232 153 1266 187
rect 1232 85 1266 119
rect 1232 17 1266 51
rect 1232 -51 1266 -17
rect 1232 -119 1266 -85
rect 1232 -187 1266 -153
rect 1232 -255 1266 -221
rect 1232 -323 1266 -289
rect 1232 -391 1266 -357
rect 1232 -459 1266 -425
rect 1232 -527 1266 -493
rect 1232 -595 1266 -561
rect 1232 -663 1266 -629
rect 1232 -731 1266 -697
rect 1232 -799 1266 -765
rect 1232 -867 1266 -833
rect 1232 -935 1266 -901
rect 1232 -1003 1266 -969
rect 1232 -1071 1266 -1037
rect 1232 -1139 1266 -1105
rect 1232 -1207 1266 -1173
rect 1232 -1275 1266 -1241
rect 1232 -1343 1266 -1309
rect 1232 -1411 1266 -1377
rect 1232 -1479 1266 -1445
rect 1232 -1547 1266 -1513
rect 1232 -1615 1266 -1581
rect 1232 -1683 1266 -1649
rect 1232 -1751 1266 -1717
rect 1232 -1819 1266 -1785
rect 1232 -1887 1266 -1853
rect 1232 -1955 1266 -1921
rect 1232 -2023 1266 -1989
rect 1232 -2091 1266 -2057
rect 1232 -2159 1266 -2125
rect 1232 -2227 1266 -2193
rect 1232 -2295 1266 -2261
rect 1232 -2363 1266 -2329
rect 1232 -2431 1266 -2397
rect 1232 -2499 1266 -2465
rect 1232 -2567 1266 -2533
rect 1232 -2635 1266 -2601
rect 1232 -2703 1266 -2669
rect 1232 -2771 1266 -2737
rect 1232 -2839 1266 -2805
rect 1232 -2907 1266 -2873
rect 1232 -2975 1266 -2941
rect 1232 -3043 1266 -3009
rect 1232 -3111 1266 -3077
rect 1232 -3179 1266 -3145
rect 1232 -3247 1266 -3213
rect 1232 -3315 1266 -3281
rect 1232 -3383 1266 -3349
rect 1232 -3451 1266 -3417
rect 1232 -3519 1266 -3485
rect 1232 -3587 1266 -3553
rect 1232 -3655 1266 -3621
rect 1232 -3723 1266 -3689
rect 1232 -3791 1266 -3757
rect 1232 -3859 1266 -3825
rect 1232 -3927 1266 -3893
rect 1232 -3995 1266 -3961
rect 1232 -4063 1266 -4029
rect 1232 -4131 1266 -4097
rect 1232 -4199 1266 -4165
rect 1232 -4267 1266 -4233
rect 1232 -4335 1266 -4301
rect 1232 -4403 1266 -4369
rect 1232 -4471 1266 -4437
rect 1232 -4539 1266 -4505
rect 1232 -4607 1266 -4573
rect 1232 -4675 1266 -4641
rect 1232 -4743 1266 -4709
rect 1232 -4811 1266 -4777
rect 1232 -4879 1266 -4845
rect 1232 -4947 1266 -4913
rect 1232 -5015 1266 -4981
rect -1183 -5102 -1149 -5068
rect -1115 -5102 -1081 -5068
rect -1047 -5102 -1013 -5068
rect -979 -5102 -945 -5068
rect -651 -5102 -617 -5068
rect -583 -5102 -549 -5068
rect -515 -5102 -481 -5068
rect -447 -5102 -413 -5068
rect -119 -5102 -85 -5068
rect -51 -5102 -17 -5068
rect 17 -5102 51 -5068
rect 85 -5102 119 -5068
rect 413 -5102 447 -5068
rect 481 -5102 515 -5068
rect 549 -5102 583 -5068
rect 617 -5102 651 -5068
rect 945 -5102 979 -5068
rect 1013 -5102 1047 -5068
rect 1081 -5102 1115 -5068
rect 1149 -5102 1183 -5068
<< mvpdiode >>
rect -1164 4981 -964 5000
rect -1164 -4981 -1149 4981
rect -979 -4981 -964 4981
rect -1164 -5000 -964 -4981
rect -632 4981 -432 5000
rect -632 -4981 -617 4981
rect -447 -4981 -432 4981
rect -632 -5000 -432 -4981
rect -100 4981 100 5000
rect -100 -4981 -85 4981
rect 85 -4981 100 4981
rect -100 -5000 100 -4981
rect 432 4981 632 5000
rect 432 -4981 447 4981
rect 617 -4981 632 4981
rect 432 -5000 632 -4981
rect 964 4981 1164 5000
rect 964 -4981 979 4981
rect 1149 -4981 1164 4981
rect 964 -5000 1164 -4981
<< mvpdiodec >>
rect -1149 -4981 -979 4981
rect -617 -4981 -447 4981
rect -85 -4981 85 4981
rect 447 -4981 617 4981
rect 979 -4981 1149 4981
<< locali >>
rect -1936 5346 -1421 5740
rect 1421 5346 1936 5740
rect -1936 5295 1936 5346
rect -1936 5237 -1493 5295
rect -1542 -5237 -1493 5237
rect 1488 5237 1936 5295
rect -1330 5102 1330 5168
rect -1330 5068 -1183 5102
rect -1119 5068 -1115 5102
rect -1013 5068 -1009 5102
rect -945 5068 -651 5102
rect -587 5068 -583 5102
rect -481 5068 -477 5102
rect -413 5068 -119 5102
rect -55 5068 -51 5102
rect 51 5068 55 5102
rect 119 5068 413 5102
rect 477 5068 481 5102
rect 583 5068 587 5102
rect 651 5068 945 5102
rect 1009 5068 1013 5102
rect 1115 5068 1119 5102
rect 1183 5068 1330 5102
rect -1330 5015 -1232 5068
rect -1330 4951 -1266 5015
rect -896 5015 -700 5068
rect -1330 4947 -1232 4951
rect -1330 4845 -1266 4947
rect -1330 4841 -1232 4845
rect -1330 4777 -1266 4841
rect -1330 4769 -1232 4777
rect -1330 4709 -1266 4769
rect -1330 4697 -1232 4709
rect -1330 4641 -1266 4697
rect -1330 4625 -1232 4641
rect -1330 4573 -1266 4625
rect -1330 4553 -1232 4573
rect -1330 4505 -1266 4553
rect -1330 4481 -1232 4505
rect -1330 4437 -1266 4481
rect -1330 4409 -1232 4437
rect -1330 4369 -1266 4409
rect -1330 4337 -1232 4369
rect -1330 4301 -1266 4337
rect -1330 4267 -1232 4301
rect -1330 4231 -1266 4267
rect -1330 4199 -1232 4231
rect -1330 4159 -1266 4199
rect -1330 4131 -1232 4159
rect -1330 4087 -1266 4131
rect -1330 4063 -1232 4087
rect -1330 4015 -1266 4063
rect -1330 3995 -1232 4015
rect -1330 3943 -1266 3995
rect -1330 3927 -1232 3943
rect -1330 3871 -1266 3927
rect -1330 3859 -1232 3871
rect -1330 3799 -1266 3859
rect -1330 3791 -1232 3799
rect -1330 3727 -1266 3791
rect -1330 3723 -1232 3727
rect -1330 3621 -1266 3723
rect -1330 3617 -1232 3621
rect -1330 3553 -1266 3617
rect -1330 3545 -1232 3553
rect -1330 3485 -1266 3545
rect -1330 3473 -1232 3485
rect -1330 3417 -1266 3473
rect -1330 3401 -1232 3417
rect -1330 3349 -1266 3401
rect -1330 3329 -1232 3349
rect -1330 3281 -1266 3329
rect -1330 3257 -1232 3281
rect -1330 3213 -1266 3257
rect -1330 3185 -1232 3213
rect -1330 3145 -1266 3185
rect -1330 3113 -1232 3145
rect -1330 3077 -1266 3113
rect -1330 3043 -1232 3077
rect -1330 3007 -1266 3043
rect -1330 2975 -1232 3007
rect -1330 2935 -1266 2975
rect -1330 2907 -1232 2935
rect -1330 2863 -1266 2907
rect -1330 2839 -1232 2863
rect -1330 2791 -1266 2839
rect -1330 2771 -1232 2791
rect -1330 2719 -1266 2771
rect -1330 2703 -1232 2719
rect -1330 2647 -1266 2703
rect -1330 2635 -1232 2647
rect -1330 2575 -1266 2635
rect -1330 2567 -1232 2575
rect -1330 2503 -1266 2567
rect -1330 2499 -1232 2503
rect -1330 2397 -1266 2499
rect -1330 2393 -1232 2397
rect -1330 2329 -1266 2393
rect -1330 2321 -1232 2329
rect -1330 2261 -1266 2321
rect -1330 2249 -1232 2261
rect -1330 2193 -1266 2249
rect -1330 2177 -1232 2193
rect -1330 2125 -1266 2177
rect -1330 2105 -1232 2125
rect -1330 2057 -1266 2105
rect -1330 2033 -1232 2057
rect -1330 1989 -1266 2033
rect -1330 1961 -1232 1989
rect -1330 1921 -1266 1961
rect -1330 1889 -1232 1921
rect -1330 1853 -1266 1889
rect -1330 1819 -1232 1853
rect -1330 1783 -1266 1819
rect -1330 1751 -1232 1783
rect -1330 1711 -1266 1751
rect -1330 1683 -1232 1711
rect -1330 1639 -1266 1683
rect -1330 1615 -1232 1639
rect -1330 1567 -1266 1615
rect -1330 1547 -1232 1567
rect -1330 1495 -1266 1547
rect -1330 1479 -1232 1495
rect -1330 1423 -1266 1479
rect -1330 1411 -1232 1423
rect -1330 1351 -1266 1411
rect -1330 1343 -1232 1351
rect -1330 1279 -1266 1343
rect -1330 1275 -1232 1279
rect -1330 1173 -1266 1275
rect -1330 1169 -1232 1173
rect -1330 1105 -1266 1169
rect -1330 1097 -1232 1105
rect -1330 1037 -1266 1097
rect -1330 1025 -1232 1037
rect -1330 969 -1266 1025
rect -1330 953 -1232 969
rect -1330 901 -1266 953
rect -1330 881 -1232 901
rect -1330 833 -1266 881
rect -1330 809 -1232 833
rect -1330 765 -1266 809
rect -1330 737 -1232 765
rect -1330 697 -1266 737
rect -1330 665 -1232 697
rect -1330 629 -1266 665
rect -1330 595 -1232 629
rect -1330 559 -1266 595
rect -1330 527 -1232 559
rect -1330 487 -1266 527
rect -1330 459 -1232 487
rect -1330 415 -1266 459
rect -1330 391 -1232 415
rect -1330 343 -1266 391
rect -1330 323 -1232 343
rect -1330 271 -1266 323
rect -1330 255 -1232 271
rect -1330 199 -1266 255
rect -1330 187 -1232 199
rect -1330 127 -1266 187
rect -1330 119 -1232 127
rect -1330 55 -1266 119
rect -1330 51 -1232 55
rect -1330 -51 -1266 51
rect -1330 -55 -1232 -51
rect -1330 -119 -1266 -55
rect -1330 -127 -1232 -119
rect -1330 -187 -1266 -127
rect -1330 -199 -1232 -187
rect -1330 -255 -1266 -199
rect -1330 -271 -1232 -255
rect -1330 -323 -1266 -271
rect -1330 -343 -1232 -323
rect -1330 -391 -1266 -343
rect -1330 -415 -1232 -391
rect -1330 -459 -1266 -415
rect -1330 -487 -1232 -459
rect -1330 -527 -1266 -487
rect -1330 -559 -1232 -527
rect -1330 -595 -1266 -559
rect -1330 -629 -1232 -595
rect -1330 -665 -1266 -629
rect -1330 -697 -1232 -665
rect -1330 -737 -1266 -697
rect -1330 -765 -1232 -737
rect -1330 -809 -1266 -765
rect -1330 -833 -1232 -809
rect -1330 -881 -1266 -833
rect -1330 -901 -1232 -881
rect -1330 -953 -1266 -901
rect -1330 -969 -1232 -953
rect -1330 -1025 -1266 -969
rect -1330 -1037 -1232 -1025
rect -1330 -1097 -1266 -1037
rect -1330 -1105 -1232 -1097
rect -1330 -1169 -1266 -1105
rect -1330 -1173 -1232 -1169
rect -1330 -1275 -1266 -1173
rect -1330 -1279 -1232 -1275
rect -1330 -1343 -1266 -1279
rect -1330 -1351 -1232 -1343
rect -1330 -1411 -1266 -1351
rect -1330 -1423 -1232 -1411
rect -1330 -1479 -1266 -1423
rect -1330 -1495 -1232 -1479
rect -1330 -1547 -1266 -1495
rect -1330 -1567 -1232 -1547
rect -1330 -1615 -1266 -1567
rect -1330 -1639 -1232 -1615
rect -1330 -1683 -1266 -1639
rect -1330 -1711 -1232 -1683
rect -1330 -1751 -1266 -1711
rect -1330 -1783 -1232 -1751
rect -1330 -1819 -1266 -1783
rect -1330 -1853 -1232 -1819
rect -1330 -1889 -1266 -1853
rect -1330 -1921 -1232 -1889
rect -1330 -1961 -1266 -1921
rect -1330 -1989 -1232 -1961
rect -1330 -2033 -1266 -1989
rect -1330 -2057 -1232 -2033
rect -1330 -2105 -1266 -2057
rect -1330 -2125 -1232 -2105
rect -1330 -2177 -1266 -2125
rect -1330 -2193 -1232 -2177
rect -1330 -2249 -1266 -2193
rect -1330 -2261 -1232 -2249
rect -1330 -2321 -1266 -2261
rect -1330 -2329 -1232 -2321
rect -1330 -2393 -1266 -2329
rect -1330 -2397 -1232 -2393
rect -1330 -2499 -1266 -2397
rect -1330 -2503 -1232 -2499
rect -1330 -2567 -1266 -2503
rect -1330 -2575 -1232 -2567
rect -1330 -2635 -1266 -2575
rect -1330 -2647 -1232 -2635
rect -1330 -2703 -1266 -2647
rect -1330 -2719 -1232 -2703
rect -1330 -2771 -1266 -2719
rect -1330 -2791 -1232 -2771
rect -1330 -2839 -1266 -2791
rect -1330 -2863 -1232 -2839
rect -1330 -2907 -1266 -2863
rect -1330 -2935 -1232 -2907
rect -1330 -2975 -1266 -2935
rect -1330 -3007 -1232 -2975
rect -1330 -3043 -1266 -3007
rect -1330 -3077 -1232 -3043
rect -1330 -3113 -1266 -3077
rect -1330 -3145 -1232 -3113
rect -1330 -3185 -1266 -3145
rect -1330 -3213 -1232 -3185
rect -1330 -3257 -1266 -3213
rect -1330 -3281 -1232 -3257
rect -1330 -3329 -1266 -3281
rect -1330 -3349 -1232 -3329
rect -1330 -3401 -1266 -3349
rect -1330 -3417 -1232 -3401
rect -1330 -3473 -1266 -3417
rect -1330 -3485 -1232 -3473
rect -1330 -3545 -1266 -3485
rect -1330 -3553 -1232 -3545
rect -1330 -3617 -1266 -3553
rect -1330 -3621 -1232 -3617
rect -1330 -3723 -1266 -3621
rect -1330 -3727 -1232 -3723
rect -1330 -3791 -1266 -3727
rect -1330 -3799 -1232 -3791
rect -1330 -3859 -1266 -3799
rect -1330 -3871 -1232 -3859
rect -1330 -3927 -1266 -3871
rect -1330 -3943 -1232 -3927
rect -1330 -3995 -1266 -3943
rect -1330 -4015 -1232 -3995
rect -1330 -4063 -1266 -4015
rect -1330 -4087 -1232 -4063
rect -1330 -4131 -1266 -4087
rect -1330 -4159 -1232 -4131
rect -1330 -4199 -1266 -4159
rect -1330 -4231 -1232 -4199
rect -1330 -4267 -1266 -4231
rect -1330 -4301 -1232 -4267
rect -1330 -4337 -1266 -4301
rect -1330 -4369 -1232 -4337
rect -1330 -4409 -1266 -4369
rect -1330 -4437 -1232 -4409
rect -1330 -4481 -1266 -4437
rect -1330 -4505 -1232 -4481
rect -1330 -4553 -1266 -4505
rect -1330 -4573 -1232 -4553
rect -1330 -4625 -1266 -4573
rect -1330 -4641 -1232 -4625
rect -1330 -4697 -1266 -4641
rect -1330 -4709 -1232 -4697
rect -1330 -4769 -1266 -4709
rect -1330 -4777 -1232 -4769
rect -1330 -4841 -1266 -4777
rect -1330 -4845 -1232 -4841
rect -1330 -4947 -1266 -4845
rect -1330 -4951 -1232 -4947
rect -1330 -5015 -1266 -4951
rect -1152 4985 -976 5004
rect -1152 4981 -1117 4985
rect -1011 4981 -976 4985
rect -1152 -4981 -1149 4981
rect -979 -4981 -976 4981
rect -1152 -4985 -1117 -4981
rect -1011 -4985 -976 -4981
rect -1152 -5004 -976 -4985
rect -862 4951 -815 5015
rect -781 4951 -734 5015
rect -364 5015 -168 5068
rect -896 4947 -700 4951
rect -862 4845 -815 4947
rect -781 4845 -734 4947
rect -896 4841 -700 4845
rect -862 4777 -815 4841
rect -781 4777 -734 4841
rect -896 4769 -700 4777
rect -862 4709 -815 4769
rect -781 4709 -734 4769
rect -896 4697 -700 4709
rect -862 4641 -815 4697
rect -781 4641 -734 4697
rect -896 4625 -700 4641
rect -862 4573 -815 4625
rect -781 4573 -734 4625
rect -896 4553 -700 4573
rect -862 4505 -815 4553
rect -781 4505 -734 4553
rect -896 4481 -700 4505
rect -862 4437 -815 4481
rect -781 4437 -734 4481
rect -896 4409 -700 4437
rect -862 4369 -815 4409
rect -781 4369 -734 4409
rect -896 4337 -700 4369
rect -862 4301 -815 4337
rect -781 4301 -734 4337
rect -896 4267 -700 4301
rect -862 4231 -815 4267
rect -781 4231 -734 4267
rect -896 4199 -700 4231
rect -862 4159 -815 4199
rect -781 4159 -734 4199
rect -896 4131 -700 4159
rect -862 4087 -815 4131
rect -781 4087 -734 4131
rect -896 4063 -700 4087
rect -862 4015 -815 4063
rect -781 4015 -734 4063
rect -896 3995 -700 4015
rect -862 3943 -815 3995
rect -781 3943 -734 3995
rect -896 3927 -700 3943
rect -862 3871 -815 3927
rect -781 3871 -734 3927
rect -896 3859 -700 3871
rect -862 3799 -815 3859
rect -781 3799 -734 3859
rect -896 3791 -700 3799
rect -862 3727 -815 3791
rect -781 3727 -734 3791
rect -896 3723 -700 3727
rect -862 3621 -815 3723
rect -781 3621 -734 3723
rect -896 3617 -700 3621
rect -862 3553 -815 3617
rect -781 3553 -734 3617
rect -896 3545 -700 3553
rect -862 3485 -815 3545
rect -781 3485 -734 3545
rect -896 3473 -700 3485
rect -862 3417 -815 3473
rect -781 3417 -734 3473
rect -896 3401 -700 3417
rect -862 3349 -815 3401
rect -781 3349 -734 3401
rect -896 3329 -700 3349
rect -862 3281 -815 3329
rect -781 3281 -734 3329
rect -896 3257 -700 3281
rect -862 3213 -815 3257
rect -781 3213 -734 3257
rect -896 3185 -700 3213
rect -862 3145 -815 3185
rect -781 3145 -734 3185
rect -896 3113 -700 3145
rect -862 3077 -815 3113
rect -781 3077 -734 3113
rect -896 3043 -700 3077
rect -862 3007 -815 3043
rect -781 3007 -734 3043
rect -896 2975 -700 3007
rect -862 2935 -815 2975
rect -781 2935 -734 2975
rect -896 2907 -700 2935
rect -862 2863 -815 2907
rect -781 2863 -734 2907
rect -896 2839 -700 2863
rect -862 2791 -815 2839
rect -781 2791 -734 2839
rect -896 2771 -700 2791
rect -862 2719 -815 2771
rect -781 2719 -734 2771
rect -896 2703 -700 2719
rect -862 2647 -815 2703
rect -781 2647 -734 2703
rect -896 2635 -700 2647
rect -862 2575 -815 2635
rect -781 2575 -734 2635
rect -896 2567 -700 2575
rect -862 2503 -815 2567
rect -781 2503 -734 2567
rect -896 2499 -700 2503
rect -862 2397 -815 2499
rect -781 2397 -734 2499
rect -896 2393 -700 2397
rect -862 2329 -815 2393
rect -781 2329 -734 2393
rect -896 2321 -700 2329
rect -862 2261 -815 2321
rect -781 2261 -734 2321
rect -896 2249 -700 2261
rect -862 2193 -815 2249
rect -781 2193 -734 2249
rect -896 2177 -700 2193
rect -862 2125 -815 2177
rect -781 2125 -734 2177
rect -896 2105 -700 2125
rect -862 2057 -815 2105
rect -781 2057 -734 2105
rect -896 2033 -700 2057
rect -862 1989 -815 2033
rect -781 1989 -734 2033
rect -896 1961 -700 1989
rect -862 1921 -815 1961
rect -781 1921 -734 1961
rect -896 1889 -700 1921
rect -862 1853 -815 1889
rect -781 1853 -734 1889
rect -896 1819 -700 1853
rect -862 1783 -815 1819
rect -781 1783 -734 1819
rect -896 1751 -700 1783
rect -862 1711 -815 1751
rect -781 1711 -734 1751
rect -896 1683 -700 1711
rect -862 1639 -815 1683
rect -781 1639 -734 1683
rect -896 1615 -700 1639
rect -862 1567 -815 1615
rect -781 1567 -734 1615
rect -896 1547 -700 1567
rect -862 1495 -815 1547
rect -781 1495 -734 1547
rect -896 1479 -700 1495
rect -862 1423 -815 1479
rect -781 1423 -734 1479
rect -896 1411 -700 1423
rect -862 1351 -815 1411
rect -781 1351 -734 1411
rect -896 1343 -700 1351
rect -862 1279 -815 1343
rect -781 1279 -734 1343
rect -896 1275 -700 1279
rect -862 1173 -815 1275
rect -781 1173 -734 1275
rect -896 1169 -700 1173
rect -862 1105 -815 1169
rect -781 1105 -734 1169
rect -896 1097 -700 1105
rect -862 1037 -815 1097
rect -781 1037 -734 1097
rect -896 1025 -700 1037
rect -862 969 -815 1025
rect -781 969 -734 1025
rect -896 953 -700 969
rect -862 901 -815 953
rect -781 901 -734 953
rect -896 881 -700 901
rect -862 833 -815 881
rect -781 833 -734 881
rect -896 809 -700 833
rect -862 765 -815 809
rect -781 765 -734 809
rect -896 737 -700 765
rect -862 697 -815 737
rect -781 697 -734 737
rect -896 665 -700 697
rect -862 629 -815 665
rect -781 629 -734 665
rect -896 595 -700 629
rect -862 559 -815 595
rect -781 559 -734 595
rect -896 527 -700 559
rect -862 487 -815 527
rect -781 487 -734 527
rect -896 459 -700 487
rect -862 415 -815 459
rect -781 415 -734 459
rect -896 391 -700 415
rect -862 343 -815 391
rect -781 343 -734 391
rect -896 323 -700 343
rect -862 271 -815 323
rect -781 271 -734 323
rect -896 255 -700 271
rect -862 199 -815 255
rect -781 199 -734 255
rect -896 187 -700 199
rect -862 127 -815 187
rect -781 127 -734 187
rect -896 119 -700 127
rect -862 55 -815 119
rect -781 55 -734 119
rect -896 51 -700 55
rect -862 -51 -815 51
rect -781 -51 -734 51
rect -896 -55 -700 -51
rect -862 -119 -815 -55
rect -781 -119 -734 -55
rect -896 -127 -700 -119
rect -862 -187 -815 -127
rect -781 -187 -734 -127
rect -896 -199 -700 -187
rect -862 -255 -815 -199
rect -781 -255 -734 -199
rect -896 -271 -700 -255
rect -862 -323 -815 -271
rect -781 -323 -734 -271
rect -896 -343 -700 -323
rect -862 -391 -815 -343
rect -781 -391 -734 -343
rect -896 -415 -700 -391
rect -862 -459 -815 -415
rect -781 -459 -734 -415
rect -896 -487 -700 -459
rect -862 -527 -815 -487
rect -781 -527 -734 -487
rect -896 -559 -700 -527
rect -862 -595 -815 -559
rect -781 -595 -734 -559
rect -896 -629 -700 -595
rect -862 -665 -815 -629
rect -781 -665 -734 -629
rect -896 -697 -700 -665
rect -862 -737 -815 -697
rect -781 -737 -734 -697
rect -896 -765 -700 -737
rect -862 -809 -815 -765
rect -781 -809 -734 -765
rect -896 -833 -700 -809
rect -862 -881 -815 -833
rect -781 -881 -734 -833
rect -896 -901 -700 -881
rect -862 -953 -815 -901
rect -781 -953 -734 -901
rect -896 -969 -700 -953
rect -862 -1025 -815 -969
rect -781 -1025 -734 -969
rect -896 -1037 -700 -1025
rect -862 -1097 -815 -1037
rect -781 -1097 -734 -1037
rect -896 -1105 -700 -1097
rect -862 -1169 -815 -1105
rect -781 -1169 -734 -1105
rect -896 -1173 -700 -1169
rect -862 -1275 -815 -1173
rect -781 -1275 -734 -1173
rect -896 -1279 -700 -1275
rect -862 -1343 -815 -1279
rect -781 -1343 -734 -1279
rect -896 -1351 -700 -1343
rect -862 -1411 -815 -1351
rect -781 -1411 -734 -1351
rect -896 -1423 -700 -1411
rect -862 -1479 -815 -1423
rect -781 -1479 -734 -1423
rect -896 -1495 -700 -1479
rect -862 -1547 -815 -1495
rect -781 -1547 -734 -1495
rect -896 -1567 -700 -1547
rect -862 -1615 -815 -1567
rect -781 -1615 -734 -1567
rect -896 -1639 -700 -1615
rect -862 -1683 -815 -1639
rect -781 -1683 -734 -1639
rect -896 -1711 -700 -1683
rect -862 -1751 -815 -1711
rect -781 -1751 -734 -1711
rect -896 -1783 -700 -1751
rect -862 -1819 -815 -1783
rect -781 -1819 -734 -1783
rect -896 -1853 -700 -1819
rect -862 -1889 -815 -1853
rect -781 -1889 -734 -1853
rect -896 -1921 -700 -1889
rect -862 -1961 -815 -1921
rect -781 -1961 -734 -1921
rect -896 -1989 -700 -1961
rect -862 -2033 -815 -1989
rect -781 -2033 -734 -1989
rect -896 -2057 -700 -2033
rect -862 -2105 -815 -2057
rect -781 -2105 -734 -2057
rect -896 -2125 -700 -2105
rect -862 -2177 -815 -2125
rect -781 -2177 -734 -2125
rect -896 -2193 -700 -2177
rect -862 -2249 -815 -2193
rect -781 -2249 -734 -2193
rect -896 -2261 -700 -2249
rect -862 -2321 -815 -2261
rect -781 -2321 -734 -2261
rect -896 -2329 -700 -2321
rect -862 -2393 -815 -2329
rect -781 -2393 -734 -2329
rect -896 -2397 -700 -2393
rect -862 -2499 -815 -2397
rect -781 -2499 -734 -2397
rect -896 -2503 -700 -2499
rect -862 -2567 -815 -2503
rect -781 -2567 -734 -2503
rect -896 -2575 -700 -2567
rect -862 -2635 -815 -2575
rect -781 -2635 -734 -2575
rect -896 -2647 -700 -2635
rect -862 -2703 -815 -2647
rect -781 -2703 -734 -2647
rect -896 -2719 -700 -2703
rect -862 -2771 -815 -2719
rect -781 -2771 -734 -2719
rect -896 -2791 -700 -2771
rect -862 -2839 -815 -2791
rect -781 -2839 -734 -2791
rect -896 -2863 -700 -2839
rect -862 -2907 -815 -2863
rect -781 -2907 -734 -2863
rect -896 -2935 -700 -2907
rect -862 -2975 -815 -2935
rect -781 -2975 -734 -2935
rect -896 -3007 -700 -2975
rect -862 -3043 -815 -3007
rect -781 -3043 -734 -3007
rect -896 -3077 -700 -3043
rect -862 -3113 -815 -3077
rect -781 -3113 -734 -3077
rect -896 -3145 -700 -3113
rect -862 -3185 -815 -3145
rect -781 -3185 -734 -3145
rect -896 -3213 -700 -3185
rect -862 -3257 -815 -3213
rect -781 -3257 -734 -3213
rect -896 -3281 -700 -3257
rect -862 -3329 -815 -3281
rect -781 -3329 -734 -3281
rect -896 -3349 -700 -3329
rect -862 -3401 -815 -3349
rect -781 -3401 -734 -3349
rect -896 -3417 -700 -3401
rect -862 -3473 -815 -3417
rect -781 -3473 -734 -3417
rect -896 -3485 -700 -3473
rect -862 -3545 -815 -3485
rect -781 -3545 -734 -3485
rect -896 -3553 -700 -3545
rect -862 -3617 -815 -3553
rect -781 -3617 -734 -3553
rect -896 -3621 -700 -3617
rect -862 -3723 -815 -3621
rect -781 -3723 -734 -3621
rect -896 -3727 -700 -3723
rect -862 -3791 -815 -3727
rect -781 -3791 -734 -3727
rect -896 -3799 -700 -3791
rect -862 -3859 -815 -3799
rect -781 -3859 -734 -3799
rect -896 -3871 -700 -3859
rect -862 -3927 -815 -3871
rect -781 -3927 -734 -3871
rect -896 -3943 -700 -3927
rect -862 -3995 -815 -3943
rect -781 -3995 -734 -3943
rect -896 -4015 -700 -3995
rect -862 -4063 -815 -4015
rect -781 -4063 -734 -4015
rect -896 -4087 -700 -4063
rect -862 -4131 -815 -4087
rect -781 -4131 -734 -4087
rect -896 -4159 -700 -4131
rect -862 -4199 -815 -4159
rect -781 -4199 -734 -4159
rect -896 -4231 -700 -4199
rect -862 -4267 -815 -4231
rect -781 -4267 -734 -4231
rect -896 -4301 -700 -4267
rect -862 -4337 -815 -4301
rect -781 -4337 -734 -4301
rect -896 -4369 -700 -4337
rect -862 -4409 -815 -4369
rect -781 -4409 -734 -4369
rect -896 -4437 -700 -4409
rect -862 -4481 -815 -4437
rect -781 -4481 -734 -4437
rect -896 -4505 -700 -4481
rect -862 -4553 -815 -4505
rect -781 -4553 -734 -4505
rect -896 -4573 -700 -4553
rect -862 -4625 -815 -4573
rect -781 -4625 -734 -4573
rect -896 -4641 -700 -4625
rect -862 -4697 -815 -4641
rect -781 -4697 -734 -4641
rect -896 -4709 -700 -4697
rect -862 -4769 -815 -4709
rect -781 -4769 -734 -4709
rect -896 -4777 -700 -4769
rect -862 -4841 -815 -4777
rect -781 -4841 -734 -4777
rect -896 -4845 -700 -4841
rect -862 -4947 -815 -4845
rect -781 -4947 -734 -4845
rect -896 -4951 -700 -4947
rect -1330 -5068 -1232 -5015
rect -862 -5015 -815 -4951
rect -781 -5015 -734 -4951
rect -620 4985 -444 5004
rect -620 4981 -585 4985
rect -479 4981 -444 4985
rect -620 -4981 -617 4981
rect -447 -4981 -444 4981
rect -620 -4985 -585 -4981
rect -479 -4985 -444 -4981
rect -620 -5004 -444 -4985
rect -330 4951 -283 5015
rect -249 4951 -202 5015
rect 168 5015 364 5068
rect -364 4947 -168 4951
rect -330 4845 -283 4947
rect -249 4845 -202 4947
rect -364 4841 -168 4845
rect -330 4777 -283 4841
rect -249 4777 -202 4841
rect -364 4769 -168 4777
rect -330 4709 -283 4769
rect -249 4709 -202 4769
rect -364 4697 -168 4709
rect -330 4641 -283 4697
rect -249 4641 -202 4697
rect -364 4625 -168 4641
rect -330 4573 -283 4625
rect -249 4573 -202 4625
rect -364 4553 -168 4573
rect -330 4505 -283 4553
rect -249 4505 -202 4553
rect -364 4481 -168 4505
rect -330 4437 -283 4481
rect -249 4437 -202 4481
rect -364 4409 -168 4437
rect -330 4369 -283 4409
rect -249 4369 -202 4409
rect -364 4337 -168 4369
rect -330 4301 -283 4337
rect -249 4301 -202 4337
rect -364 4267 -168 4301
rect -330 4231 -283 4267
rect -249 4231 -202 4267
rect -364 4199 -168 4231
rect -330 4159 -283 4199
rect -249 4159 -202 4199
rect -364 4131 -168 4159
rect -330 4087 -283 4131
rect -249 4087 -202 4131
rect -364 4063 -168 4087
rect -330 4015 -283 4063
rect -249 4015 -202 4063
rect -364 3995 -168 4015
rect -330 3943 -283 3995
rect -249 3943 -202 3995
rect -364 3927 -168 3943
rect -330 3871 -283 3927
rect -249 3871 -202 3927
rect -364 3859 -168 3871
rect -330 3799 -283 3859
rect -249 3799 -202 3859
rect -364 3791 -168 3799
rect -330 3727 -283 3791
rect -249 3727 -202 3791
rect -364 3723 -168 3727
rect -330 3621 -283 3723
rect -249 3621 -202 3723
rect -364 3617 -168 3621
rect -330 3553 -283 3617
rect -249 3553 -202 3617
rect -364 3545 -168 3553
rect -330 3485 -283 3545
rect -249 3485 -202 3545
rect -364 3473 -168 3485
rect -330 3417 -283 3473
rect -249 3417 -202 3473
rect -364 3401 -168 3417
rect -330 3349 -283 3401
rect -249 3349 -202 3401
rect -364 3329 -168 3349
rect -330 3281 -283 3329
rect -249 3281 -202 3329
rect -364 3257 -168 3281
rect -330 3213 -283 3257
rect -249 3213 -202 3257
rect -364 3185 -168 3213
rect -330 3145 -283 3185
rect -249 3145 -202 3185
rect -364 3113 -168 3145
rect -330 3077 -283 3113
rect -249 3077 -202 3113
rect -364 3043 -168 3077
rect -330 3007 -283 3043
rect -249 3007 -202 3043
rect -364 2975 -168 3007
rect -330 2935 -283 2975
rect -249 2935 -202 2975
rect -364 2907 -168 2935
rect -330 2863 -283 2907
rect -249 2863 -202 2907
rect -364 2839 -168 2863
rect -330 2791 -283 2839
rect -249 2791 -202 2839
rect -364 2771 -168 2791
rect -330 2719 -283 2771
rect -249 2719 -202 2771
rect -364 2703 -168 2719
rect -330 2647 -283 2703
rect -249 2647 -202 2703
rect -364 2635 -168 2647
rect -330 2575 -283 2635
rect -249 2575 -202 2635
rect -364 2567 -168 2575
rect -330 2503 -283 2567
rect -249 2503 -202 2567
rect -364 2499 -168 2503
rect -330 2397 -283 2499
rect -249 2397 -202 2499
rect -364 2393 -168 2397
rect -330 2329 -283 2393
rect -249 2329 -202 2393
rect -364 2321 -168 2329
rect -330 2261 -283 2321
rect -249 2261 -202 2321
rect -364 2249 -168 2261
rect -330 2193 -283 2249
rect -249 2193 -202 2249
rect -364 2177 -168 2193
rect -330 2125 -283 2177
rect -249 2125 -202 2177
rect -364 2105 -168 2125
rect -330 2057 -283 2105
rect -249 2057 -202 2105
rect -364 2033 -168 2057
rect -330 1989 -283 2033
rect -249 1989 -202 2033
rect -364 1961 -168 1989
rect -330 1921 -283 1961
rect -249 1921 -202 1961
rect -364 1889 -168 1921
rect -330 1853 -283 1889
rect -249 1853 -202 1889
rect -364 1819 -168 1853
rect -330 1783 -283 1819
rect -249 1783 -202 1819
rect -364 1751 -168 1783
rect -330 1711 -283 1751
rect -249 1711 -202 1751
rect -364 1683 -168 1711
rect -330 1639 -283 1683
rect -249 1639 -202 1683
rect -364 1615 -168 1639
rect -330 1567 -283 1615
rect -249 1567 -202 1615
rect -364 1547 -168 1567
rect -330 1495 -283 1547
rect -249 1495 -202 1547
rect -364 1479 -168 1495
rect -330 1423 -283 1479
rect -249 1423 -202 1479
rect -364 1411 -168 1423
rect -330 1351 -283 1411
rect -249 1351 -202 1411
rect -364 1343 -168 1351
rect -330 1279 -283 1343
rect -249 1279 -202 1343
rect -364 1275 -168 1279
rect -330 1173 -283 1275
rect -249 1173 -202 1275
rect -364 1169 -168 1173
rect -330 1105 -283 1169
rect -249 1105 -202 1169
rect -364 1097 -168 1105
rect -330 1037 -283 1097
rect -249 1037 -202 1097
rect -364 1025 -168 1037
rect -330 969 -283 1025
rect -249 969 -202 1025
rect -364 953 -168 969
rect -330 901 -283 953
rect -249 901 -202 953
rect -364 881 -168 901
rect -330 833 -283 881
rect -249 833 -202 881
rect -364 809 -168 833
rect -330 765 -283 809
rect -249 765 -202 809
rect -364 737 -168 765
rect -330 697 -283 737
rect -249 697 -202 737
rect -364 665 -168 697
rect -330 629 -283 665
rect -249 629 -202 665
rect -364 595 -168 629
rect -330 559 -283 595
rect -249 559 -202 595
rect -364 527 -168 559
rect -330 487 -283 527
rect -249 487 -202 527
rect -364 459 -168 487
rect -330 415 -283 459
rect -249 415 -202 459
rect -364 391 -168 415
rect -330 343 -283 391
rect -249 343 -202 391
rect -364 323 -168 343
rect -330 271 -283 323
rect -249 271 -202 323
rect -364 255 -168 271
rect -330 199 -283 255
rect -249 199 -202 255
rect -364 187 -168 199
rect -330 127 -283 187
rect -249 127 -202 187
rect -364 119 -168 127
rect -330 55 -283 119
rect -249 55 -202 119
rect -364 51 -168 55
rect -330 -51 -283 51
rect -249 -51 -202 51
rect -364 -55 -168 -51
rect -330 -119 -283 -55
rect -249 -119 -202 -55
rect -364 -127 -168 -119
rect -330 -187 -283 -127
rect -249 -187 -202 -127
rect -364 -199 -168 -187
rect -330 -255 -283 -199
rect -249 -255 -202 -199
rect -364 -271 -168 -255
rect -330 -323 -283 -271
rect -249 -323 -202 -271
rect -364 -343 -168 -323
rect -330 -391 -283 -343
rect -249 -391 -202 -343
rect -364 -415 -168 -391
rect -330 -459 -283 -415
rect -249 -459 -202 -415
rect -364 -487 -168 -459
rect -330 -527 -283 -487
rect -249 -527 -202 -487
rect -364 -559 -168 -527
rect -330 -595 -283 -559
rect -249 -595 -202 -559
rect -364 -629 -168 -595
rect -330 -665 -283 -629
rect -249 -665 -202 -629
rect -364 -697 -168 -665
rect -330 -737 -283 -697
rect -249 -737 -202 -697
rect -364 -765 -168 -737
rect -330 -809 -283 -765
rect -249 -809 -202 -765
rect -364 -833 -168 -809
rect -330 -881 -283 -833
rect -249 -881 -202 -833
rect -364 -901 -168 -881
rect -330 -953 -283 -901
rect -249 -953 -202 -901
rect -364 -969 -168 -953
rect -330 -1025 -283 -969
rect -249 -1025 -202 -969
rect -364 -1037 -168 -1025
rect -330 -1097 -283 -1037
rect -249 -1097 -202 -1037
rect -364 -1105 -168 -1097
rect -330 -1169 -283 -1105
rect -249 -1169 -202 -1105
rect -364 -1173 -168 -1169
rect -330 -1275 -283 -1173
rect -249 -1275 -202 -1173
rect -364 -1279 -168 -1275
rect -330 -1343 -283 -1279
rect -249 -1343 -202 -1279
rect -364 -1351 -168 -1343
rect -330 -1411 -283 -1351
rect -249 -1411 -202 -1351
rect -364 -1423 -168 -1411
rect -330 -1479 -283 -1423
rect -249 -1479 -202 -1423
rect -364 -1495 -168 -1479
rect -330 -1547 -283 -1495
rect -249 -1547 -202 -1495
rect -364 -1567 -168 -1547
rect -330 -1615 -283 -1567
rect -249 -1615 -202 -1567
rect -364 -1639 -168 -1615
rect -330 -1683 -283 -1639
rect -249 -1683 -202 -1639
rect -364 -1711 -168 -1683
rect -330 -1751 -283 -1711
rect -249 -1751 -202 -1711
rect -364 -1783 -168 -1751
rect -330 -1819 -283 -1783
rect -249 -1819 -202 -1783
rect -364 -1853 -168 -1819
rect -330 -1889 -283 -1853
rect -249 -1889 -202 -1853
rect -364 -1921 -168 -1889
rect -330 -1961 -283 -1921
rect -249 -1961 -202 -1921
rect -364 -1989 -168 -1961
rect -330 -2033 -283 -1989
rect -249 -2033 -202 -1989
rect -364 -2057 -168 -2033
rect -330 -2105 -283 -2057
rect -249 -2105 -202 -2057
rect -364 -2125 -168 -2105
rect -330 -2177 -283 -2125
rect -249 -2177 -202 -2125
rect -364 -2193 -168 -2177
rect -330 -2249 -283 -2193
rect -249 -2249 -202 -2193
rect -364 -2261 -168 -2249
rect -330 -2321 -283 -2261
rect -249 -2321 -202 -2261
rect -364 -2329 -168 -2321
rect -330 -2393 -283 -2329
rect -249 -2393 -202 -2329
rect -364 -2397 -168 -2393
rect -330 -2499 -283 -2397
rect -249 -2499 -202 -2397
rect -364 -2503 -168 -2499
rect -330 -2567 -283 -2503
rect -249 -2567 -202 -2503
rect -364 -2575 -168 -2567
rect -330 -2635 -283 -2575
rect -249 -2635 -202 -2575
rect -364 -2647 -168 -2635
rect -330 -2703 -283 -2647
rect -249 -2703 -202 -2647
rect -364 -2719 -168 -2703
rect -330 -2771 -283 -2719
rect -249 -2771 -202 -2719
rect -364 -2791 -168 -2771
rect -330 -2839 -283 -2791
rect -249 -2839 -202 -2791
rect -364 -2863 -168 -2839
rect -330 -2907 -283 -2863
rect -249 -2907 -202 -2863
rect -364 -2935 -168 -2907
rect -330 -2975 -283 -2935
rect -249 -2975 -202 -2935
rect -364 -3007 -168 -2975
rect -330 -3043 -283 -3007
rect -249 -3043 -202 -3007
rect -364 -3077 -168 -3043
rect -330 -3113 -283 -3077
rect -249 -3113 -202 -3077
rect -364 -3145 -168 -3113
rect -330 -3185 -283 -3145
rect -249 -3185 -202 -3145
rect -364 -3213 -168 -3185
rect -330 -3257 -283 -3213
rect -249 -3257 -202 -3213
rect -364 -3281 -168 -3257
rect -330 -3329 -283 -3281
rect -249 -3329 -202 -3281
rect -364 -3349 -168 -3329
rect -330 -3401 -283 -3349
rect -249 -3401 -202 -3349
rect -364 -3417 -168 -3401
rect -330 -3473 -283 -3417
rect -249 -3473 -202 -3417
rect -364 -3485 -168 -3473
rect -330 -3545 -283 -3485
rect -249 -3545 -202 -3485
rect -364 -3553 -168 -3545
rect -330 -3617 -283 -3553
rect -249 -3617 -202 -3553
rect -364 -3621 -168 -3617
rect -330 -3723 -283 -3621
rect -249 -3723 -202 -3621
rect -364 -3727 -168 -3723
rect -330 -3791 -283 -3727
rect -249 -3791 -202 -3727
rect -364 -3799 -168 -3791
rect -330 -3859 -283 -3799
rect -249 -3859 -202 -3799
rect -364 -3871 -168 -3859
rect -330 -3927 -283 -3871
rect -249 -3927 -202 -3871
rect -364 -3943 -168 -3927
rect -330 -3995 -283 -3943
rect -249 -3995 -202 -3943
rect -364 -4015 -168 -3995
rect -330 -4063 -283 -4015
rect -249 -4063 -202 -4015
rect -364 -4087 -168 -4063
rect -330 -4131 -283 -4087
rect -249 -4131 -202 -4087
rect -364 -4159 -168 -4131
rect -330 -4199 -283 -4159
rect -249 -4199 -202 -4159
rect -364 -4231 -168 -4199
rect -330 -4267 -283 -4231
rect -249 -4267 -202 -4231
rect -364 -4301 -168 -4267
rect -330 -4337 -283 -4301
rect -249 -4337 -202 -4301
rect -364 -4369 -168 -4337
rect -330 -4409 -283 -4369
rect -249 -4409 -202 -4369
rect -364 -4437 -168 -4409
rect -330 -4481 -283 -4437
rect -249 -4481 -202 -4437
rect -364 -4505 -168 -4481
rect -330 -4553 -283 -4505
rect -249 -4553 -202 -4505
rect -364 -4573 -168 -4553
rect -330 -4625 -283 -4573
rect -249 -4625 -202 -4573
rect -364 -4641 -168 -4625
rect -330 -4697 -283 -4641
rect -249 -4697 -202 -4641
rect -364 -4709 -168 -4697
rect -330 -4769 -283 -4709
rect -249 -4769 -202 -4709
rect -364 -4777 -168 -4769
rect -330 -4841 -283 -4777
rect -249 -4841 -202 -4777
rect -364 -4845 -168 -4841
rect -330 -4947 -283 -4845
rect -249 -4947 -202 -4845
rect -364 -4951 -168 -4947
rect -896 -5068 -700 -5015
rect -330 -5015 -283 -4951
rect -249 -5015 -202 -4951
rect -88 4985 88 5004
rect -88 4981 -53 4985
rect 53 4981 88 4985
rect -88 -4981 -85 4981
rect 85 -4981 88 4981
rect -88 -4985 -53 -4981
rect 53 -4985 88 -4981
rect -88 -5004 88 -4985
rect 202 4951 249 5015
rect 283 4951 330 5015
rect 700 5015 896 5068
rect 168 4947 364 4951
rect 202 4845 249 4947
rect 283 4845 330 4947
rect 168 4841 364 4845
rect 202 4777 249 4841
rect 283 4777 330 4841
rect 168 4769 364 4777
rect 202 4709 249 4769
rect 283 4709 330 4769
rect 168 4697 364 4709
rect 202 4641 249 4697
rect 283 4641 330 4697
rect 168 4625 364 4641
rect 202 4573 249 4625
rect 283 4573 330 4625
rect 168 4553 364 4573
rect 202 4505 249 4553
rect 283 4505 330 4553
rect 168 4481 364 4505
rect 202 4437 249 4481
rect 283 4437 330 4481
rect 168 4409 364 4437
rect 202 4369 249 4409
rect 283 4369 330 4409
rect 168 4337 364 4369
rect 202 4301 249 4337
rect 283 4301 330 4337
rect 168 4267 364 4301
rect 202 4231 249 4267
rect 283 4231 330 4267
rect 168 4199 364 4231
rect 202 4159 249 4199
rect 283 4159 330 4199
rect 168 4131 364 4159
rect 202 4087 249 4131
rect 283 4087 330 4131
rect 168 4063 364 4087
rect 202 4015 249 4063
rect 283 4015 330 4063
rect 168 3995 364 4015
rect 202 3943 249 3995
rect 283 3943 330 3995
rect 168 3927 364 3943
rect 202 3871 249 3927
rect 283 3871 330 3927
rect 168 3859 364 3871
rect 202 3799 249 3859
rect 283 3799 330 3859
rect 168 3791 364 3799
rect 202 3727 249 3791
rect 283 3727 330 3791
rect 168 3723 364 3727
rect 202 3621 249 3723
rect 283 3621 330 3723
rect 168 3617 364 3621
rect 202 3553 249 3617
rect 283 3553 330 3617
rect 168 3545 364 3553
rect 202 3485 249 3545
rect 283 3485 330 3545
rect 168 3473 364 3485
rect 202 3417 249 3473
rect 283 3417 330 3473
rect 168 3401 364 3417
rect 202 3349 249 3401
rect 283 3349 330 3401
rect 168 3329 364 3349
rect 202 3281 249 3329
rect 283 3281 330 3329
rect 168 3257 364 3281
rect 202 3213 249 3257
rect 283 3213 330 3257
rect 168 3185 364 3213
rect 202 3145 249 3185
rect 283 3145 330 3185
rect 168 3113 364 3145
rect 202 3077 249 3113
rect 283 3077 330 3113
rect 168 3043 364 3077
rect 202 3007 249 3043
rect 283 3007 330 3043
rect 168 2975 364 3007
rect 202 2935 249 2975
rect 283 2935 330 2975
rect 168 2907 364 2935
rect 202 2863 249 2907
rect 283 2863 330 2907
rect 168 2839 364 2863
rect 202 2791 249 2839
rect 283 2791 330 2839
rect 168 2771 364 2791
rect 202 2719 249 2771
rect 283 2719 330 2771
rect 168 2703 364 2719
rect 202 2647 249 2703
rect 283 2647 330 2703
rect 168 2635 364 2647
rect 202 2575 249 2635
rect 283 2575 330 2635
rect 168 2567 364 2575
rect 202 2503 249 2567
rect 283 2503 330 2567
rect 168 2499 364 2503
rect 202 2397 249 2499
rect 283 2397 330 2499
rect 168 2393 364 2397
rect 202 2329 249 2393
rect 283 2329 330 2393
rect 168 2321 364 2329
rect 202 2261 249 2321
rect 283 2261 330 2321
rect 168 2249 364 2261
rect 202 2193 249 2249
rect 283 2193 330 2249
rect 168 2177 364 2193
rect 202 2125 249 2177
rect 283 2125 330 2177
rect 168 2105 364 2125
rect 202 2057 249 2105
rect 283 2057 330 2105
rect 168 2033 364 2057
rect 202 1989 249 2033
rect 283 1989 330 2033
rect 168 1961 364 1989
rect 202 1921 249 1961
rect 283 1921 330 1961
rect 168 1889 364 1921
rect 202 1853 249 1889
rect 283 1853 330 1889
rect 168 1819 364 1853
rect 202 1783 249 1819
rect 283 1783 330 1819
rect 168 1751 364 1783
rect 202 1711 249 1751
rect 283 1711 330 1751
rect 168 1683 364 1711
rect 202 1639 249 1683
rect 283 1639 330 1683
rect 168 1615 364 1639
rect 202 1567 249 1615
rect 283 1567 330 1615
rect 168 1547 364 1567
rect 202 1495 249 1547
rect 283 1495 330 1547
rect 168 1479 364 1495
rect 202 1423 249 1479
rect 283 1423 330 1479
rect 168 1411 364 1423
rect 202 1351 249 1411
rect 283 1351 330 1411
rect 168 1343 364 1351
rect 202 1279 249 1343
rect 283 1279 330 1343
rect 168 1275 364 1279
rect 202 1173 249 1275
rect 283 1173 330 1275
rect 168 1169 364 1173
rect 202 1105 249 1169
rect 283 1105 330 1169
rect 168 1097 364 1105
rect 202 1037 249 1097
rect 283 1037 330 1097
rect 168 1025 364 1037
rect 202 969 249 1025
rect 283 969 330 1025
rect 168 953 364 969
rect 202 901 249 953
rect 283 901 330 953
rect 168 881 364 901
rect 202 833 249 881
rect 283 833 330 881
rect 168 809 364 833
rect 202 765 249 809
rect 283 765 330 809
rect 168 737 364 765
rect 202 697 249 737
rect 283 697 330 737
rect 168 665 364 697
rect 202 629 249 665
rect 283 629 330 665
rect 168 595 364 629
rect 202 559 249 595
rect 283 559 330 595
rect 168 527 364 559
rect 202 487 249 527
rect 283 487 330 527
rect 168 459 364 487
rect 202 415 249 459
rect 283 415 330 459
rect 168 391 364 415
rect 202 343 249 391
rect 283 343 330 391
rect 168 323 364 343
rect 202 271 249 323
rect 283 271 330 323
rect 168 255 364 271
rect 202 199 249 255
rect 283 199 330 255
rect 168 187 364 199
rect 202 127 249 187
rect 283 127 330 187
rect 168 119 364 127
rect 202 55 249 119
rect 283 55 330 119
rect 168 51 364 55
rect 202 -51 249 51
rect 283 -51 330 51
rect 168 -55 364 -51
rect 202 -119 249 -55
rect 283 -119 330 -55
rect 168 -127 364 -119
rect 202 -187 249 -127
rect 283 -187 330 -127
rect 168 -199 364 -187
rect 202 -255 249 -199
rect 283 -255 330 -199
rect 168 -271 364 -255
rect 202 -323 249 -271
rect 283 -323 330 -271
rect 168 -343 364 -323
rect 202 -391 249 -343
rect 283 -391 330 -343
rect 168 -415 364 -391
rect 202 -459 249 -415
rect 283 -459 330 -415
rect 168 -487 364 -459
rect 202 -527 249 -487
rect 283 -527 330 -487
rect 168 -559 364 -527
rect 202 -595 249 -559
rect 283 -595 330 -559
rect 168 -629 364 -595
rect 202 -665 249 -629
rect 283 -665 330 -629
rect 168 -697 364 -665
rect 202 -737 249 -697
rect 283 -737 330 -697
rect 168 -765 364 -737
rect 202 -809 249 -765
rect 283 -809 330 -765
rect 168 -833 364 -809
rect 202 -881 249 -833
rect 283 -881 330 -833
rect 168 -901 364 -881
rect 202 -953 249 -901
rect 283 -953 330 -901
rect 168 -969 364 -953
rect 202 -1025 249 -969
rect 283 -1025 330 -969
rect 168 -1037 364 -1025
rect 202 -1097 249 -1037
rect 283 -1097 330 -1037
rect 168 -1105 364 -1097
rect 202 -1169 249 -1105
rect 283 -1169 330 -1105
rect 168 -1173 364 -1169
rect 202 -1275 249 -1173
rect 283 -1275 330 -1173
rect 168 -1279 364 -1275
rect 202 -1343 249 -1279
rect 283 -1343 330 -1279
rect 168 -1351 364 -1343
rect 202 -1411 249 -1351
rect 283 -1411 330 -1351
rect 168 -1423 364 -1411
rect 202 -1479 249 -1423
rect 283 -1479 330 -1423
rect 168 -1495 364 -1479
rect 202 -1547 249 -1495
rect 283 -1547 330 -1495
rect 168 -1567 364 -1547
rect 202 -1615 249 -1567
rect 283 -1615 330 -1567
rect 168 -1639 364 -1615
rect 202 -1683 249 -1639
rect 283 -1683 330 -1639
rect 168 -1711 364 -1683
rect 202 -1751 249 -1711
rect 283 -1751 330 -1711
rect 168 -1783 364 -1751
rect 202 -1819 249 -1783
rect 283 -1819 330 -1783
rect 168 -1853 364 -1819
rect 202 -1889 249 -1853
rect 283 -1889 330 -1853
rect 168 -1921 364 -1889
rect 202 -1961 249 -1921
rect 283 -1961 330 -1921
rect 168 -1989 364 -1961
rect 202 -2033 249 -1989
rect 283 -2033 330 -1989
rect 168 -2057 364 -2033
rect 202 -2105 249 -2057
rect 283 -2105 330 -2057
rect 168 -2125 364 -2105
rect 202 -2177 249 -2125
rect 283 -2177 330 -2125
rect 168 -2193 364 -2177
rect 202 -2249 249 -2193
rect 283 -2249 330 -2193
rect 168 -2261 364 -2249
rect 202 -2321 249 -2261
rect 283 -2321 330 -2261
rect 168 -2329 364 -2321
rect 202 -2393 249 -2329
rect 283 -2393 330 -2329
rect 168 -2397 364 -2393
rect 202 -2499 249 -2397
rect 283 -2499 330 -2397
rect 168 -2503 364 -2499
rect 202 -2567 249 -2503
rect 283 -2567 330 -2503
rect 168 -2575 364 -2567
rect 202 -2635 249 -2575
rect 283 -2635 330 -2575
rect 168 -2647 364 -2635
rect 202 -2703 249 -2647
rect 283 -2703 330 -2647
rect 168 -2719 364 -2703
rect 202 -2771 249 -2719
rect 283 -2771 330 -2719
rect 168 -2791 364 -2771
rect 202 -2839 249 -2791
rect 283 -2839 330 -2791
rect 168 -2863 364 -2839
rect 202 -2907 249 -2863
rect 283 -2907 330 -2863
rect 168 -2935 364 -2907
rect 202 -2975 249 -2935
rect 283 -2975 330 -2935
rect 168 -3007 364 -2975
rect 202 -3043 249 -3007
rect 283 -3043 330 -3007
rect 168 -3077 364 -3043
rect 202 -3113 249 -3077
rect 283 -3113 330 -3077
rect 168 -3145 364 -3113
rect 202 -3185 249 -3145
rect 283 -3185 330 -3145
rect 168 -3213 364 -3185
rect 202 -3257 249 -3213
rect 283 -3257 330 -3213
rect 168 -3281 364 -3257
rect 202 -3329 249 -3281
rect 283 -3329 330 -3281
rect 168 -3349 364 -3329
rect 202 -3401 249 -3349
rect 283 -3401 330 -3349
rect 168 -3417 364 -3401
rect 202 -3473 249 -3417
rect 283 -3473 330 -3417
rect 168 -3485 364 -3473
rect 202 -3545 249 -3485
rect 283 -3545 330 -3485
rect 168 -3553 364 -3545
rect 202 -3617 249 -3553
rect 283 -3617 330 -3553
rect 168 -3621 364 -3617
rect 202 -3723 249 -3621
rect 283 -3723 330 -3621
rect 168 -3727 364 -3723
rect 202 -3791 249 -3727
rect 283 -3791 330 -3727
rect 168 -3799 364 -3791
rect 202 -3859 249 -3799
rect 283 -3859 330 -3799
rect 168 -3871 364 -3859
rect 202 -3927 249 -3871
rect 283 -3927 330 -3871
rect 168 -3943 364 -3927
rect 202 -3995 249 -3943
rect 283 -3995 330 -3943
rect 168 -4015 364 -3995
rect 202 -4063 249 -4015
rect 283 -4063 330 -4015
rect 168 -4087 364 -4063
rect 202 -4131 249 -4087
rect 283 -4131 330 -4087
rect 168 -4159 364 -4131
rect 202 -4199 249 -4159
rect 283 -4199 330 -4159
rect 168 -4231 364 -4199
rect 202 -4267 249 -4231
rect 283 -4267 330 -4231
rect 168 -4301 364 -4267
rect 202 -4337 249 -4301
rect 283 -4337 330 -4301
rect 168 -4369 364 -4337
rect 202 -4409 249 -4369
rect 283 -4409 330 -4369
rect 168 -4437 364 -4409
rect 202 -4481 249 -4437
rect 283 -4481 330 -4437
rect 168 -4505 364 -4481
rect 202 -4553 249 -4505
rect 283 -4553 330 -4505
rect 168 -4573 364 -4553
rect 202 -4625 249 -4573
rect 283 -4625 330 -4573
rect 168 -4641 364 -4625
rect 202 -4697 249 -4641
rect 283 -4697 330 -4641
rect 168 -4709 364 -4697
rect 202 -4769 249 -4709
rect 283 -4769 330 -4709
rect 168 -4777 364 -4769
rect 202 -4841 249 -4777
rect 283 -4841 330 -4777
rect 168 -4845 364 -4841
rect 202 -4947 249 -4845
rect 283 -4947 330 -4845
rect 168 -4951 364 -4947
rect -364 -5068 -168 -5015
rect 202 -5015 249 -4951
rect 283 -5015 330 -4951
rect 444 4985 620 5004
rect 444 4981 479 4985
rect 585 4981 620 4985
rect 444 -4981 447 4981
rect 617 -4981 620 4981
rect 444 -4985 479 -4981
rect 585 -4985 620 -4981
rect 444 -5004 620 -4985
rect 734 4951 781 5015
rect 815 4951 862 5015
rect 1232 5015 1330 5068
rect 700 4947 896 4951
rect 734 4845 781 4947
rect 815 4845 862 4947
rect 700 4841 896 4845
rect 734 4777 781 4841
rect 815 4777 862 4841
rect 700 4769 896 4777
rect 734 4709 781 4769
rect 815 4709 862 4769
rect 700 4697 896 4709
rect 734 4641 781 4697
rect 815 4641 862 4697
rect 700 4625 896 4641
rect 734 4573 781 4625
rect 815 4573 862 4625
rect 700 4553 896 4573
rect 734 4505 781 4553
rect 815 4505 862 4553
rect 700 4481 896 4505
rect 734 4437 781 4481
rect 815 4437 862 4481
rect 700 4409 896 4437
rect 734 4369 781 4409
rect 815 4369 862 4409
rect 700 4337 896 4369
rect 734 4301 781 4337
rect 815 4301 862 4337
rect 700 4267 896 4301
rect 734 4231 781 4267
rect 815 4231 862 4267
rect 700 4199 896 4231
rect 734 4159 781 4199
rect 815 4159 862 4199
rect 700 4131 896 4159
rect 734 4087 781 4131
rect 815 4087 862 4131
rect 700 4063 896 4087
rect 734 4015 781 4063
rect 815 4015 862 4063
rect 700 3995 896 4015
rect 734 3943 781 3995
rect 815 3943 862 3995
rect 700 3927 896 3943
rect 734 3871 781 3927
rect 815 3871 862 3927
rect 700 3859 896 3871
rect 734 3799 781 3859
rect 815 3799 862 3859
rect 700 3791 896 3799
rect 734 3727 781 3791
rect 815 3727 862 3791
rect 700 3723 896 3727
rect 734 3621 781 3723
rect 815 3621 862 3723
rect 700 3617 896 3621
rect 734 3553 781 3617
rect 815 3553 862 3617
rect 700 3545 896 3553
rect 734 3485 781 3545
rect 815 3485 862 3545
rect 700 3473 896 3485
rect 734 3417 781 3473
rect 815 3417 862 3473
rect 700 3401 896 3417
rect 734 3349 781 3401
rect 815 3349 862 3401
rect 700 3329 896 3349
rect 734 3281 781 3329
rect 815 3281 862 3329
rect 700 3257 896 3281
rect 734 3213 781 3257
rect 815 3213 862 3257
rect 700 3185 896 3213
rect 734 3145 781 3185
rect 815 3145 862 3185
rect 700 3113 896 3145
rect 734 3077 781 3113
rect 815 3077 862 3113
rect 700 3043 896 3077
rect 734 3007 781 3043
rect 815 3007 862 3043
rect 700 2975 896 3007
rect 734 2935 781 2975
rect 815 2935 862 2975
rect 700 2907 896 2935
rect 734 2863 781 2907
rect 815 2863 862 2907
rect 700 2839 896 2863
rect 734 2791 781 2839
rect 815 2791 862 2839
rect 700 2771 896 2791
rect 734 2719 781 2771
rect 815 2719 862 2771
rect 700 2703 896 2719
rect 734 2647 781 2703
rect 815 2647 862 2703
rect 700 2635 896 2647
rect 734 2575 781 2635
rect 815 2575 862 2635
rect 700 2567 896 2575
rect 734 2503 781 2567
rect 815 2503 862 2567
rect 700 2499 896 2503
rect 734 2397 781 2499
rect 815 2397 862 2499
rect 700 2393 896 2397
rect 734 2329 781 2393
rect 815 2329 862 2393
rect 700 2321 896 2329
rect 734 2261 781 2321
rect 815 2261 862 2321
rect 700 2249 896 2261
rect 734 2193 781 2249
rect 815 2193 862 2249
rect 700 2177 896 2193
rect 734 2125 781 2177
rect 815 2125 862 2177
rect 700 2105 896 2125
rect 734 2057 781 2105
rect 815 2057 862 2105
rect 700 2033 896 2057
rect 734 1989 781 2033
rect 815 1989 862 2033
rect 700 1961 896 1989
rect 734 1921 781 1961
rect 815 1921 862 1961
rect 700 1889 896 1921
rect 734 1853 781 1889
rect 815 1853 862 1889
rect 700 1819 896 1853
rect 734 1783 781 1819
rect 815 1783 862 1819
rect 700 1751 896 1783
rect 734 1711 781 1751
rect 815 1711 862 1751
rect 700 1683 896 1711
rect 734 1639 781 1683
rect 815 1639 862 1683
rect 700 1615 896 1639
rect 734 1567 781 1615
rect 815 1567 862 1615
rect 700 1547 896 1567
rect 734 1495 781 1547
rect 815 1495 862 1547
rect 700 1479 896 1495
rect 734 1423 781 1479
rect 815 1423 862 1479
rect 700 1411 896 1423
rect 734 1351 781 1411
rect 815 1351 862 1411
rect 700 1343 896 1351
rect 734 1279 781 1343
rect 815 1279 862 1343
rect 700 1275 896 1279
rect 734 1173 781 1275
rect 815 1173 862 1275
rect 700 1169 896 1173
rect 734 1105 781 1169
rect 815 1105 862 1169
rect 700 1097 896 1105
rect 734 1037 781 1097
rect 815 1037 862 1097
rect 700 1025 896 1037
rect 734 969 781 1025
rect 815 969 862 1025
rect 700 953 896 969
rect 734 901 781 953
rect 815 901 862 953
rect 700 881 896 901
rect 734 833 781 881
rect 815 833 862 881
rect 700 809 896 833
rect 734 765 781 809
rect 815 765 862 809
rect 700 737 896 765
rect 734 697 781 737
rect 815 697 862 737
rect 700 665 896 697
rect 734 629 781 665
rect 815 629 862 665
rect 700 595 896 629
rect 734 559 781 595
rect 815 559 862 595
rect 700 527 896 559
rect 734 487 781 527
rect 815 487 862 527
rect 700 459 896 487
rect 734 415 781 459
rect 815 415 862 459
rect 700 391 896 415
rect 734 343 781 391
rect 815 343 862 391
rect 700 323 896 343
rect 734 271 781 323
rect 815 271 862 323
rect 700 255 896 271
rect 734 199 781 255
rect 815 199 862 255
rect 700 187 896 199
rect 734 127 781 187
rect 815 127 862 187
rect 700 119 896 127
rect 734 55 781 119
rect 815 55 862 119
rect 700 51 896 55
rect 734 -51 781 51
rect 815 -51 862 51
rect 700 -55 896 -51
rect 734 -119 781 -55
rect 815 -119 862 -55
rect 700 -127 896 -119
rect 734 -187 781 -127
rect 815 -187 862 -127
rect 700 -199 896 -187
rect 734 -255 781 -199
rect 815 -255 862 -199
rect 700 -271 896 -255
rect 734 -323 781 -271
rect 815 -323 862 -271
rect 700 -343 896 -323
rect 734 -391 781 -343
rect 815 -391 862 -343
rect 700 -415 896 -391
rect 734 -459 781 -415
rect 815 -459 862 -415
rect 700 -487 896 -459
rect 734 -527 781 -487
rect 815 -527 862 -487
rect 700 -559 896 -527
rect 734 -595 781 -559
rect 815 -595 862 -559
rect 700 -629 896 -595
rect 734 -665 781 -629
rect 815 -665 862 -629
rect 700 -697 896 -665
rect 734 -737 781 -697
rect 815 -737 862 -697
rect 700 -765 896 -737
rect 734 -809 781 -765
rect 815 -809 862 -765
rect 700 -833 896 -809
rect 734 -881 781 -833
rect 815 -881 862 -833
rect 700 -901 896 -881
rect 734 -953 781 -901
rect 815 -953 862 -901
rect 700 -969 896 -953
rect 734 -1025 781 -969
rect 815 -1025 862 -969
rect 700 -1037 896 -1025
rect 734 -1097 781 -1037
rect 815 -1097 862 -1037
rect 700 -1105 896 -1097
rect 734 -1169 781 -1105
rect 815 -1169 862 -1105
rect 700 -1173 896 -1169
rect 734 -1275 781 -1173
rect 815 -1275 862 -1173
rect 700 -1279 896 -1275
rect 734 -1343 781 -1279
rect 815 -1343 862 -1279
rect 700 -1351 896 -1343
rect 734 -1411 781 -1351
rect 815 -1411 862 -1351
rect 700 -1423 896 -1411
rect 734 -1479 781 -1423
rect 815 -1479 862 -1423
rect 700 -1495 896 -1479
rect 734 -1547 781 -1495
rect 815 -1547 862 -1495
rect 700 -1567 896 -1547
rect 734 -1615 781 -1567
rect 815 -1615 862 -1567
rect 700 -1639 896 -1615
rect 734 -1683 781 -1639
rect 815 -1683 862 -1639
rect 700 -1711 896 -1683
rect 734 -1751 781 -1711
rect 815 -1751 862 -1711
rect 700 -1783 896 -1751
rect 734 -1819 781 -1783
rect 815 -1819 862 -1783
rect 700 -1853 896 -1819
rect 734 -1889 781 -1853
rect 815 -1889 862 -1853
rect 700 -1921 896 -1889
rect 734 -1961 781 -1921
rect 815 -1961 862 -1921
rect 700 -1989 896 -1961
rect 734 -2033 781 -1989
rect 815 -2033 862 -1989
rect 700 -2057 896 -2033
rect 734 -2105 781 -2057
rect 815 -2105 862 -2057
rect 700 -2125 896 -2105
rect 734 -2177 781 -2125
rect 815 -2177 862 -2125
rect 700 -2193 896 -2177
rect 734 -2249 781 -2193
rect 815 -2249 862 -2193
rect 700 -2261 896 -2249
rect 734 -2321 781 -2261
rect 815 -2321 862 -2261
rect 700 -2329 896 -2321
rect 734 -2393 781 -2329
rect 815 -2393 862 -2329
rect 700 -2397 896 -2393
rect 734 -2499 781 -2397
rect 815 -2499 862 -2397
rect 700 -2503 896 -2499
rect 734 -2567 781 -2503
rect 815 -2567 862 -2503
rect 700 -2575 896 -2567
rect 734 -2635 781 -2575
rect 815 -2635 862 -2575
rect 700 -2647 896 -2635
rect 734 -2703 781 -2647
rect 815 -2703 862 -2647
rect 700 -2719 896 -2703
rect 734 -2771 781 -2719
rect 815 -2771 862 -2719
rect 700 -2791 896 -2771
rect 734 -2839 781 -2791
rect 815 -2839 862 -2791
rect 700 -2863 896 -2839
rect 734 -2907 781 -2863
rect 815 -2907 862 -2863
rect 700 -2935 896 -2907
rect 734 -2975 781 -2935
rect 815 -2975 862 -2935
rect 700 -3007 896 -2975
rect 734 -3043 781 -3007
rect 815 -3043 862 -3007
rect 700 -3077 896 -3043
rect 734 -3113 781 -3077
rect 815 -3113 862 -3077
rect 700 -3145 896 -3113
rect 734 -3185 781 -3145
rect 815 -3185 862 -3145
rect 700 -3213 896 -3185
rect 734 -3257 781 -3213
rect 815 -3257 862 -3213
rect 700 -3281 896 -3257
rect 734 -3329 781 -3281
rect 815 -3329 862 -3281
rect 700 -3349 896 -3329
rect 734 -3401 781 -3349
rect 815 -3401 862 -3349
rect 700 -3417 896 -3401
rect 734 -3473 781 -3417
rect 815 -3473 862 -3417
rect 700 -3485 896 -3473
rect 734 -3545 781 -3485
rect 815 -3545 862 -3485
rect 700 -3553 896 -3545
rect 734 -3617 781 -3553
rect 815 -3617 862 -3553
rect 700 -3621 896 -3617
rect 734 -3723 781 -3621
rect 815 -3723 862 -3621
rect 700 -3727 896 -3723
rect 734 -3791 781 -3727
rect 815 -3791 862 -3727
rect 700 -3799 896 -3791
rect 734 -3859 781 -3799
rect 815 -3859 862 -3799
rect 700 -3871 896 -3859
rect 734 -3927 781 -3871
rect 815 -3927 862 -3871
rect 700 -3943 896 -3927
rect 734 -3995 781 -3943
rect 815 -3995 862 -3943
rect 700 -4015 896 -3995
rect 734 -4063 781 -4015
rect 815 -4063 862 -4015
rect 700 -4087 896 -4063
rect 734 -4131 781 -4087
rect 815 -4131 862 -4087
rect 700 -4159 896 -4131
rect 734 -4199 781 -4159
rect 815 -4199 862 -4159
rect 700 -4231 896 -4199
rect 734 -4267 781 -4231
rect 815 -4267 862 -4231
rect 700 -4301 896 -4267
rect 734 -4337 781 -4301
rect 815 -4337 862 -4301
rect 700 -4369 896 -4337
rect 734 -4409 781 -4369
rect 815 -4409 862 -4369
rect 700 -4437 896 -4409
rect 734 -4481 781 -4437
rect 815 -4481 862 -4437
rect 700 -4505 896 -4481
rect 734 -4553 781 -4505
rect 815 -4553 862 -4505
rect 700 -4573 896 -4553
rect 734 -4625 781 -4573
rect 815 -4625 862 -4573
rect 700 -4641 896 -4625
rect 734 -4697 781 -4641
rect 815 -4697 862 -4641
rect 700 -4709 896 -4697
rect 734 -4769 781 -4709
rect 815 -4769 862 -4709
rect 700 -4777 896 -4769
rect 734 -4841 781 -4777
rect 815 -4841 862 -4777
rect 700 -4845 896 -4841
rect 734 -4947 781 -4845
rect 815 -4947 862 -4845
rect 700 -4951 896 -4947
rect 168 -5068 364 -5015
rect 734 -5015 781 -4951
rect 815 -5015 862 -4951
rect 976 4985 1152 5004
rect 976 4981 1011 4985
rect 1117 4981 1152 4985
rect 976 -4981 979 4981
rect 1149 -4981 1152 4981
rect 976 -4985 1011 -4981
rect 1117 -4985 1152 -4981
rect 976 -5004 1152 -4985
rect 1266 4951 1330 5015
rect 1232 4947 1330 4951
rect 1266 4845 1330 4947
rect 1232 4841 1330 4845
rect 1266 4777 1330 4841
rect 1232 4769 1330 4777
rect 1266 4709 1330 4769
rect 1232 4697 1330 4709
rect 1266 4641 1330 4697
rect 1232 4625 1330 4641
rect 1266 4573 1330 4625
rect 1232 4553 1330 4573
rect 1266 4505 1330 4553
rect 1232 4481 1330 4505
rect 1266 4437 1330 4481
rect 1232 4409 1330 4437
rect 1266 4369 1330 4409
rect 1232 4337 1330 4369
rect 1266 4301 1330 4337
rect 1232 4267 1330 4301
rect 1266 4231 1330 4267
rect 1232 4199 1330 4231
rect 1266 4159 1330 4199
rect 1232 4131 1330 4159
rect 1266 4087 1330 4131
rect 1232 4063 1330 4087
rect 1266 4015 1330 4063
rect 1232 3995 1330 4015
rect 1266 3943 1330 3995
rect 1232 3927 1330 3943
rect 1266 3871 1330 3927
rect 1232 3859 1330 3871
rect 1266 3799 1330 3859
rect 1232 3791 1330 3799
rect 1266 3727 1330 3791
rect 1232 3723 1330 3727
rect 1266 3621 1330 3723
rect 1232 3617 1330 3621
rect 1266 3553 1330 3617
rect 1232 3545 1330 3553
rect 1266 3485 1330 3545
rect 1232 3473 1330 3485
rect 1266 3417 1330 3473
rect 1232 3401 1330 3417
rect 1266 3349 1330 3401
rect 1232 3329 1330 3349
rect 1266 3281 1330 3329
rect 1232 3257 1330 3281
rect 1266 3213 1330 3257
rect 1232 3185 1330 3213
rect 1266 3145 1330 3185
rect 1232 3113 1330 3145
rect 1266 3077 1330 3113
rect 1232 3043 1330 3077
rect 1266 3007 1330 3043
rect 1232 2975 1330 3007
rect 1266 2935 1330 2975
rect 1232 2907 1330 2935
rect 1266 2863 1330 2907
rect 1232 2839 1330 2863
rect 1266 2791 1330 2839
rect 1232 2771 1330 2791
rect 1266 2719 1330 2771
rect 1232 2703 1330 2719
rect 1266 2647 1330 2703
rect 1232 2635 1330 2647
rect 1266 2575 1330 2635
rect 1232 2567 1330 2575
rect 1266 2503 1330 2567
rect 1232 2499 1330 2503
rect 1266 2397 1330 2499
rect 1232 2393 1330 2397
rect 1266 2329 1330 2393
rect 1232 2321 1330 2329
rect 1266 2261 1330 2321
rect 1232 2249 1330 2261
rect 1266 2193 1330 2249
rect 1232 2177 1330 2193
rect 1266 2125 1330 2177
rect 1232 2105 1330 2125
rect 1266 2057 1330 2105
rect 1232 2033 1330 2057
rect 1266 1989 1330 2033
rect 1232 1961 1330 1989
rect 1266 1921 1330 1961
rect 1232 1889 1330 1921
rect 1266 1853 1330 1889
rect 1232 1819 1330 1853
rect 1266 1783 1330 1819
rect 1232 1751 1330 1783
rect 1266 1711 1330 1751
rect 1232 1683 1330 1711
rect 1266 1639 1330 1683
rect 1232 1615 1330 1639
rect 1266 1567 1330 1615
rect 1232 1547 1330 1567
rect 1266 1495 1330 1547
rect 1232 1479 1330 1495
rect 1266 1423 1330 1479
rect 1232 1411 1330 1423
rect 1266 1351 1330 1411
rect 1232 1343 1330 1351
rect 1266 1279 1330 1343
rect 1232 1275 1330 1279
rect 1266 1173 1330 1275
rect 1232 1169 1330 1173
rect 1266 1105 1330 1169
rect 1232 1097 1330 1105
rect 1266 1037 1330 1097
rect 1232 1025 1330 1037
rect 1266 969 1330 1025
rect 1232 953 1330 969
rect 1266 901 1330 953
rect 1232 881 1330 901
rect 1266 833 1330 881
rect 1232 809 1330 833
rect 1266 765 1330 809
rect 1232 737 1330 765
rect 1266 697 1330 737
rect 1232 665 1330 697
rect 1266 629 1330 665
rect 1232 595 1330 629
rect 1266 559 1330 595
rect 1232 527 1330 559
rect 1266 487 1330 527
rect 1232 459 1330 487
rect 1266 415 1330 459
rect 1232 391 1330 415
rect 1266 343 1330 391
rect 1232 323 1330 343
rect 1266 271 1330 323
rect 1232 255 1330 271
rect 1266 199 1330 255
rect 1232 187 1330 199
rect 1266 127 1330 187
rect 1232 119 1330 127
rect 1266 55 1330 119
rect 1232 51 1330 55
rect 1266 -51 1330 51
rect 1232 -55 1330 -51
rect 1266 -119 1330 -55
rect 1232 -127 1330 -119
rect 1266 -187 1330 -127
rect 1232 -199 1330 -187
rect 1266 -255 1330 -199
rect 1232 -271 1330 -255
rect 1266 -323 1330 -271
rect 1232 -343 1330 -323
rect 1266 -391 1330 -343
rect 1232 -415 1330 -391
rect 1266 -459 1330 -415
rect 1232 -487 1330 -459
rect 1266 -527 1330 -487
rect 1232 -559 1330 -527
rect 1266 -595 1330 -559
rect 1232 -629 1330 -595
rect 1266 -665 1330 -629
rect 1232 -697 1330 -665
rect 1266 -737 1330 -697
rect 1232 -765 1330 -737
rect 1266 -809 1330 -765
rect 1232 -833 1330 -809
rect 1266 -881 1330 -833
rect 1232 -901 1330 -881
rect 1266 -953 1330 -901
rect 1232 -969 1330 -953
rect 1266 -1025 1330 -969
rect 1232 -1037 1330 -1025
rect 1266 -1097 1330 -1037
rect 1232 -1105 1330 -1097
rect 1266 -1169 1330 -1105
rect 1232 -1173 1330 -1169
rect 1266 -1275 1330 -1173
rect 1232 -1279 1330 -1275
rect 1266 -1343 1330 -1279
rect 1232 -1351 1330 -1343
rect 1266 -1411 1330 -1351
rect 1232 -1423 1330 -1411
rect 1266 -1479 1330 -1423
rect 1232 -1495 1330 -1479
rect 1266 -1547 1330 -1495
rect 1232 -1567 1330 -1547
rect 1266 -1615 1330 -1567
rect 1232 -1639 1330 -1615
rect 1266 -1683 1330 -1639
rect 1232 -1711 1330 -1683
rect 1266 -1751 1330 -1711
rect 1232 -1783 1330 -1751
rect 1266 -1819 1330 -1783
rect 1232 -1853 1330 -1819
rect 1266 -1889 1330 -1853
rect 1232 -1921 1330 -1889
rect 1266 -1961 1330 -1921
rect 1232 -1989 1330 -1961
rect 1266 -2033 1330 -1989
rect 1232 -2057 1330 -2033
rect 1266 -2105 1330 -2057
rect 1232 -2125 1330 -2105
rect 1266 -2177 1330 -2125
rect 1232 -2193 1330 -2177
rect 1266 -2249 1330 -2193
rect 1232 -2261 1330 -2249
rect 1266 -2321 1330 -2261
rect 1232 -2329 1330 -2321
rect 1266 -2393 1330 -2329
rect 1232 -2397 1330 -2393
rect 1266 -2499 1330 -2397
rect 1232 -2503 1330 -2499
rect 1266 -2567 1330 -2503
rect 1232 -2575 1330 -2567
rect 1266 -2635 1330 -2575
rect 1232 -2647 1330 -2635
rect 1266 -2703 1330 -2647
rect 1232 -2719 1330 -2703
rect 1266 -2771 1330 -2719
rect 1232 -2791 1330 -2771
rect 1266 -2839 1330 -2791
rect 1232 -2863 1330 -2839
rect 1266 -2907 1330 -2863
rect 1232 -2935 1330 -2907
rect 1266 -2975 1330 -2935
rect 1232 -3007 1330 -2975
rect 1266 -3043 1330 -3007
rect 1232 -3077 1330 -3043
rect 1266 -3113 1330 -3077
rect 1232 -3145 1330 -3113
rect 1266 -3185 1330 -3145
rect 1232 -3213 1330 -3185
rect 1266 -3257 1330 -3213
rect 1232 -3281 1330 -3257
rect 1266 -3329 1330 -3281
rect 1232 -3349 1330 -3329
rect 1266 -3401 1330 -3349
rect 1232 -3417 1330 -3401
rect 1266 -3473 1330 -3417
rect 1232 -3485 1330 -3473
rect 1266 -3545 1330 -3485
rect 1232 -3553 1330 -3545
rect 1266 -3617 1330 -3553
rect 1232 -3621 1330 -3617
rect 1266 -3723 1330 -3621
rect 1232 -3727 1330 -3723
rect 1266 -3791 1330 -3727
rect 1232 -3799 1330 -3791
rect 1266 -3859 1330 -3799
rect 1232 -3871 1330 -3859
rect 1266 -3927 1330 -3871
rect 1232 -3943 1330 -3927
rect 1266 -3995 1330 -3943
rect 1232 -4015 1330 -3995
rect 1266 -4063 1330 -4015
rect 1232 -4087 1330 -4063
rect 1266 -4131 1330 -4087
rect 1232 -4159 1330 -4131
rect 1266 -4199 1330 -4159
rect 1232 -4231 1330 -4199
rect 1266 -4267 1330 -4231
rect 1232 -4301 1330 -4267
rect 1266 -4337 1330 -4301
rect 1232 -4369 1330 -4337
rect 1266 -4409 1330 -4369
rect 1232 -4437 1330 -4409
rect 1266 -4481 1330 -4437
rect 1232 -4505 1330 -4481
rect 1266 -4553 1330 -4505
rect 1232 -4573 1330 -4553
rect 1266 -4625 1330 -4573
rect 1232 -4641 1330 -4625
rect 1266 -4697 1330 -4641
rect 1232 -4709 1330 -4697
rect 1266 -4769 1330 -4709
rect 1232 -4777 1330 -4769
rect 1266 -4841 1330 -4777
rect 1232 -4845 1330 -4841
rect 1266 -4947 1330 -4845
rect 1232 -4951 1330 -4947
rect 700 -5068 896 -5015
rect 1266 -5015 1330 -4951
rect 1232 -5068 1330 -5015
rect -1330 -5102 -1183 -5068
rect -1119 -5102 -1115 -5068
rect -1013 -5102 -1009 -5068
rect -945 -5102 -651 -5068
rect -587 -5102 -583 -5068
rect -481 -5102 -477 -5068
rect -413 -5102 -119 -5068
rect -55 -5102 -51 -5068
rect 51 -5102 55 -5068
rect 119 -5102 413 -5068
rect 477 -5102 481 -5068
rect 583 -5102 587 -5068
rect 651 -5102 945 -5068
rect 1009 -5102 1013 -5068
rect 1115 -5102 1119 -5068
rect 1183 -5102 1330 -5068
rect -1330 -5168 1330 -5102
rect -1936 -5286 -1493 -5237
rect 1488 -5237 1542 5237
rect 1488 -5286 1936 -5237
rect -1936 -5346 1936 -5286
rect -1936 -5740 -1421 -5346
rect 1421 -5740 1936 -5346
<< viali >>
rect -1421 5730 1421 5740
rect -1421 5356 -1411 5730
rect -1411 5356 1411 5730
rect 1411 5356 1421 5730
rect -1421 5346 1421 5356
rect -1936 5219 -1542 5237
rect -1936 -5219 -1926 5219
rect -1926 -5219 -1552 5219
rect -1552 -5219 -1542 5219
rect -1936 -5237 -1542 -5219
rect -1153 5068 -1149 5102
rect -1149 5068 -1119 5102
rect -1081 5068 -1047 5102
rect -1009 5068 -979 5102
rect -979 5068 -975 5102
rect -621 5068 -617 5102
rect -617 5068 -587 5102
rect -549 5068 -515 5102
rect -477 5068 -447 5102
rect -447 5068 -443 5102
rect -89 5068 -85 5102
rect -85 5068 -55 5102
rect -17 5068 17 5102
rect 55 5068 85 5102
rect 85 5068 89 5102
rect 443 5068 447 5102
rect 447 5068 477 5102
rect 515 5068 549 5102
rect 587 5068 617 5102
rect 617 5068 621 5102
rect 975 5068 979 5102
rect 979 5068 1009 5102
rect 1047 5068 1081 5102
rect 1119 5068 1149 5102
rect 1149 5068 1153 5102
rect -1266 4981 -1232 4985
rect -1266 4951 -1232 4981
rect -1266 4879 -1232 4913
rect -1266 4811 -1232 4841
rect -1266 4807 -1232 4811
rect -1266 4743 -1232 4769
rect -1266 4735 -1232 4743
rect -1266 4675 -1232 4697
rect -1266 4663 -1232 4675
rect -1266 4607 -1232 4625
rect -1266 4591 -1232 4607
rect -1266 4539 -1232 4553
rect -1266 4519 -1232 4539
rect -1266 4471 -1232 4481
rect -1266 4447 -1232 4471
rect -1266 4403 -1232 4409
rect -1266 4375 -1232 4403
rect -1266 4335 -1232 4337
rect -1266 4303 -1232 4335
rect -1266 4233 -1232 4265
rect -1266 4231 -1232 4233
rect -1266 4165 -1232 4193
rect -1266 4159 -1232 4165
rect -1266 4097 -1232 4121
rect -1266 4087 -1232 4097
rect -1266 4029 -1232 4049
rect -1266 4015 -1232 4029
rect -1266 3961 -1232 3977
rect -1266 3943 -1232 3961
rect -1266 3893 -1232 3905
rect -1266 3871 -1232 3893
rect -1266 3825 -1232 3833
rect -1266 3799 -1232 3825
rect -1266 3757 -1232 3761
rect -1266 3727 -1232 3757
rect -1266 3655 -1232 3689
rect -1266 3587 -1232 3617
rect -1266 3583 -1232 3587
rect -1266 3519 -1232 3545
rect -1266 3511 -1232 3519
rect -1266 3451 -1232 3473
rect -1266 3439 -1232 3451
rect -1266 3383 -1232 3401
rect -1266 3367 -1232 3383
rect -1266 3315 -1232 3329
rect -1266 3295 -1232 3315
rect -1266 3247 -1232 3257
rect -1266 3223 -1232 3247
rect -1266 3179 -1232 3185
rect -1266 3151 -1232 3179
rect -1266 3111 -1232 3113
rect -1266 3079 -1232 3111
rect -1266 3009 -1232 3041
rect -1266 3007 -1232 3009
rect -1266 2941 -1232 2969
rect -1266 2935 -1232 2941
rect -1266 2873 -1232 2897
rect -1266 2863 -1232 2873
rect -1266 2805 -1232 2825
rect -1266 2791 -1232 2805
rect -1266 2737 -1232 2753
rect -1266 2719 -1232 2737
rect -1266 2669 -1232 2681
rect -1266 2647 -1232 2669
rect -1266 2601 -1232 2609
rect -1266 2575 -1232 2601
rect -1266 2533 -1232 2537
rect -1266 2503 -1232 2533
rect -1266 2431 -1232 2465
rect -1266 2363 -1232 2393
rect -1266 2359 -1232 2363
rect -1266 2295 -1232 2321
rect -1266 2287 -1232 2295
rect -1266 2227 -1232 2249
rect -1266 2215 -1232 2227
rect -1266 2159 -1232 2177
rect -1266 2143 -1232 2159
rect -1266 2091 -1232 2105
rect -1266 2071 -1232 2091
rect -1266 2023 -1232 2033
rect -1266 1999 -1232 2023
rect -1266 1955 -1232 1961
rect -1266 1927 -1232 1955
rect -1266 1887 -1232 1889
rect -1266 1855 -1232 1887
rect -1266 1785 -1232 1817
rect -1266 1783 -1232 1785
rect -1266 1717 -1232 1745
rect -1266 1711 -1232 1717
rect -1266 1649 -1232 1673
rect -1266 1639 -1232 1649
rect -1266 1581 -1232 1601
rect -1266 1567 -1232 1581
rect -1266 1513 -1232 1529
rect -1266 1495 -1232 1513
rect -1266 1445 -1232 1457
rect -1266 1423 -1232 1445
rect -1266 1377 -1232 1385
rect -1266 1351 -1232 1377
rect -1266 1309 -1232 1313
rect -1266 1279 -1232 1309
rect -1266 1207 -1232 1241
rect -1266 1139 -1232 1169
rect -1266 1135 -1232 1139
rect -1266 1071 -1232 1097
rect -1266 1063 -1232 1071
rect -1266 1003 -1232 1025
rect -1266 991 -1232 1003
rect -1266 935 -1232 953
rect -1266 919 -1232 935
rect -1266 867 -1232 881
rect -1266 847 -1232 867
rect -1266 799 -1232 809
rect -1266 775 -1232 799
rect -1266 731 -1232 737
rect -1266 703 -1232 731
rect -1266 663 -1232 665
rect -1266 631 -1232 663
rect -1266 561 -1232 593
rect -1266 559 -1232 561
rect -1266 493 -1232 521
rect -1266 487 -1232 493
rect -1266 425 -1232 449
rect -1266 415 -1232 425
rect -1266 357 -1232 377
rect -1266 343 -1232 357
rect -1266 289 -1232 305
rect -1266 271 -1232 289
rect -1266 221 -1232 233
rect -1266 199 -1232 221
rect -1266 153 -1232 161
rect -1266 127 -1232 153
rect -1266 85 -1232 89
rect -1266 55 -1232 85
rect -1266 -17 -1232 17
rect -1266 -85 -1232 -55
rect -1266 -89 -1232 -85
rect -1266 -153 -1232 -127
rect -1266 -161 -1232 -153
rect -1266 -221 -1232 -199
rect -1266 -233 -1232 -221
rect -1266 -289 -1232 -271
rect -1266 -305 -1232 -289
rect -1266 -357 -1232 -343
rect -1266 -377 -1232 -357
rect -1266 -425 -1232 -415
rect -1266 -449 -1232 -425
rect -1266 -493 -1232 -487
rect -1266 -521 -1232 -493
rect -1266 -561 -1232 -559
rect -1266 -593 -1232 -561
rect -1266 -663 -1232 -631
rect -1266 -665 -1232 -663
rect -1266 -731 -1232 -703
rect -1266 -737 -1232 -731
rect -1266 -799 -1232 -775
rect -1266 -809 -1232 -799
rect -1266 -867 -1232 -847
rect -1266 -881 -1232 -867
rect -1266 -935 -1232 -919
rect -1266 -953 -1232 -935
rect -1266 -1003 -1232 -991
rect -1266 -1025 -1232 -1003
rect -1266 -1071 -1232 -1063
rect -1266 -1097 -1232 -1071
rect -1266 -1139 -1232 -1135
rect -1266 -1169 -1232 -1139
rect -1266 -1241 -1232 -1207
rect -1266 -1309 -1232 -1279
rect -1266 -1313 -1232 -1309
rect -1266 -1377 -1232 -1351
rect -1266 -1385 -1232 -1377
rect -1266 -1445 -1232 -1423
rect -1266 -1457 -1232 -1445
rect -1266 -1513 -1232 -1495
rect -1266 -1529 -1232 -1513
rect -1266 -1581 -1232 -1567
rect -1266 -1601 -1232 -1581
rect -1266 -1649 -1232 -1639
rect -1266 -1673 -1232 -1649
rect -1266 -1717 -1232 -1711
rect -1266 -1745 -1232 -1717
rect -1266 -1785 -1232 -1783
rect -1266 -1817 -1232 -1785
rect -1266 -1887 -1232 -1855
rect -1266 -1889 -1232 -1887
rect -1266 -1955 -1232 -1927
rect -1266 -1961 -1232 -1955
rect -1266 -2023 -1232 -1999
rect -1266 -2033 -1232 -2023
rect -1266 -2091 -1232 -2071
rect -1266 -2105 -1232 -2091
rect -1266 -2159 -1232 -2143
rect -1266 -2177 -1232 -2159
rect -1266 -2227 -1232 -2215
rect -1266 -2249 -1232 -2227
rect -1266 -2295 -1232 -2287
rect -1266 -2321 -1232 -2295
rect -1266 -2363 -1232 -2359
rect -1266 -2393 -1232 -2363
rect -1266 -2465 -1232 -2431
rect -1266 -2533 -1232 -2503
rect -1266 -2537 -1232 -2533
rect -1266 -2601 -1232 -2575
rect -1266 -2609 -1232 -2601
rect -1266 -2669 -1232 -2647
rect -1266 -2681 -1232 -2669
rect -1266 -2737 -1232 -2719
rect -1266 -2753 -1232 -2737
rect -1266 -2805 -1232 -2791
rect -1266 -2825 -1232 -2805
rect -1266 -2873 -1232 -2863
rect -1266 -2897 -1232 -2873
rect -1266 -2941 -1232 -2935
rect -1266 -2969 -1232 -2941
rect -1266 -3009 -1232 -3007
rect -1266 -3041 -1232 -3009
rect -1266 -3111 -1232 -3079
rect -1266 -3113 -1232 -3111
rect -1266 -3179 -1232 -3151
rect -1266 -3185 -1232 -3179
rect -1266 -3247 -1232 -3223
rect -1266 -3257 -1232 -3247
rect -1266 -3315 -1232 -3295
rect -1266 -3329 -1232 -3315
rect -1266 -3383 -1232 -3367
rect -1266 -3401 -1232 -3383
rect -1266 -3451 -1232 -3439
rect -1266 -3473 -1232 -3451
rect -1266 -3519 -1232 -3511
rect -1266 -3545 -1232 -3519
rect -1266 -3587 -1232 -3583
rect -1266 -3617 -1232 -3587
rect -1266 -3689 -1232 -3655
rect -1266 -3757 -1232 -3727
rect -1266 -3761 -1232 -3757
rect -1266 -3825 -1232 -3799
rect -1266 -3833 -1232 -3825
rect -1266 -3893 -1232 -3871
rect -1266 -3905 -1232 -3893
rect -1266 -3961 -1232 -3943
rect -1266 -3977 -1232 -3961
rect -1266 -4029 -1232 -4015
rect -1266 -4049 -1232 -4029
rect -1266 -4097 -1232 -4087
rect -1266 -4121 -1232 -4097
rect -1266 -4165 -1232 -4159
rect -1266 -4193 -1232 -4165
rect -1266 -4233 -1232 -4231
rect -1266 -4265 -1232 -4233
rect -1266 -4335 -1232 -4303
rect -1266 -4337 -1232 -4335
rect -1266 -4403 -1232 -4375
rect -1266 -4409 -1232 -4403
rect -1266 -4471 -1232 -4447
rect -1266 -4481 -1232 -4471
rect -1266 -4539 -1232 -4519
rect -1266 -4553 -1232 -4539
rect -1266 -4607 -1232 -4591
rect -1266 -4625 -1232 -4607
rect -1266 -4675 -1232 -4663
rect -1266 -4697 -1232 -4675
rect -1266 -4743 -1232 -4735
rect -1266 -4769 -1232 -4743
rect -1266 -4811 -1232 -4807
rect -1266 -4841 -1232 -4811
rect -1266 -4913 -1232 -4879
rect -1266 -4981 -1232 -4951
rect -1266 -4985 -1232 -4981
rect -1117 4981 -1011 4985
rect -1117 -4981 -1011 4981
rect -1117 -4985 -1011 -4981
rect -896 4981 -862 4985
rect -896 4951 -862 4981
rect -815 4981 -781 4985
rect -815 4951 -781 4981
rect -734 4981 -700 4985
rect -734 4951 -700 4981
rect -896 4879 -862 4913
rect -815 4879 -781 4913
rect -734 4879 -700 4913
rect -896 4811 -862 4841
rect -896 4807 -862 4811
rect -815 4811 -781 4841
rect -815 4807 -781 4811
rect -734 4811 -700 4841
rect -734 4807 -700 4811
rect -896 4743 -862 4769
rect -896 4735 -862 4743
rect -815 4743 -781 4769
rect -815 4735 -781 4743
rect -734 4743 -700 4769
rect -734 4735 -700 4743
rect -896 4675 -862 4697
rect -896 4663 -862 4675
rect -815 4675 -781 4697
rect -815 4663 -781 4675
rect -734 4675 -700 4697
rect -734 4663 -700 4675
rect -896 4607 -862 4625
rect -896 4591 -862 4607
rect -815 4607 -781 4625
rect -815 4591 -781 4607
rect -734 4607 -700 4625
rect -734 4591 -700 4607
rect -896 4539 -862 4553
rect -896 4519 -862 4539
rect -815 4539 -781 4553
rect -815 4519 -781 4539
rect -734 4539 -700 4553
rect -734 4519 -700 4539
rect -896 4471 -862 4481
rect -896 4447 -862 4471
rect -815 4471 -781 4481
rect -815 4447 -781 4471
rect -734 4471 -700 4481
rect -734 4447 -700 4471
rect -896 4403 -862 4409
rect -896 4375 -862 4403
rect -815 4403 -781 4409
rect -815 4375 -781 4403
rect -734 4403 -700 4409
rect -734 4375 -700 4403
rect -896 4335 -862 4337
rect -896 4303 -862 4335
rect -815 4335 -781 4337
rect -815 4303 -781 4335
rect -734 4335 -700 4337
rect -734 4303 -700 4335
rect -896 4233 -862 4265
rect -896 4231 -862 4233
rect -815 4233 -781 4265
rect -815 4231 -781 4233
rect -734 4233 -700 4265
rect -734 4231 -700 4233
rect -896 4165 -862 4193
rect -896 4159 -862 4165
rect -815 4165 -781 4193
rect -815 4159 -781 4165
rect -734 4165 -700 4193
rect -734 4159 -700 4165
rect -896 4097 -862 4121
rect -896 4087 -862 4097
rect -815 4097 -781 4121
rect -815 4087 -781 4097
rect -734 4097 -700 4121
rect -734 4087 -700 4097
rect -896 4029 -862 4049
rect -896 4015 -862 4029
rect -815 4029 -781 4049
rect -815 4015 -781 4029
rect -734 4029 -700 4049
rect -734 4015 -700 4029
rect -896 3961 -862 3977
rect -896 3943 -862 3961
rect -815 3961 -781 3977
rect -815 3943 -781 3961
rect -734 3961 -700 3977
rect -734 3943 -700 3961
rect -896 3893 -862 3905
rect -896 3871 -862 3893
rect -815 3893 -781 3905
rect -815 3871 -781 3893
rect -734 3893 -700 3905
rect -734 3871 -700 3893
rect -896 3825 -862 3833
rect -896 3799 -862 3825
rect -815 3825 -781 3833
rect -815 3799 -781 3825
rect -734 3825 -700 3833
rect -734 3799 -700 3825
rect -896 3757 -862 3761
rect -896 3727 -862 3757
rect -815 3757 -781 3761
rect -815 3727 -781 3757
rect -734 3757 -700 3761
rect -734 3727 -700 3757
rect -896 3655 -862 3689
rect -815 3655 -781 3689
rect -734 3655 -700 3689
rect -896 3587 -862 3617
rect -896 3583 -862 3587
rect -815 3587 -781 3617
rect -815 3583 -781 3587
rect -734 3587 -700 3617
rect -734 3583 -700 3587
rect -896 3519 -862 3545
rect -896 3511 -862 3519
rect -815 3519 -781 3545
rect -815 3511 -781 3519
rect -734 3519 -700 3545
rect -734 3511 -700 3519
rect -896 3451 -862 3473
rect -896 3439 -862 3451
rect -815 3451 -781 3473
rect -815 3439 -781 3451
rect -734 3451 -700 3473
rect -734 3439 -700 3451
rect -896 3383 -862 3401
rect -896 3367 -862 3383
rect -815 3383 -781 3401
rect -815 3367 -781 3383
rect -734 3383 -700 3401
rect -734 3367 -700 3383
rect -896 3315 -862 3329
rect -896 3295 -862 3315
rect -815 3315 -781 3329
rect -815 3295 -781 3315
rect -734 3315 -700 3329
rect -734 3295 -700 3315
rect -896 3247 -862 3257
rect -896 3223 -862 3247
rect -815 3247 -781 3257
rect -815 3223 -781 3247
rect -734 3247 -700 3257
rect -734 3223 -700 3247
rect -896 3179 -862 3185
rect -896 3151 -862 3179
rect -815 3179 -781 3185
rect -815 3151 -781 3179
rect -734 3179 -700 3185
rect -734 3151 -700 3179
rect -896 3111 -862 3113
rect -896 3079 -862 3111
rect -815 3111 -781 3113
rect -815 3079 -781 3111
rect -734 3111 -700 3113
rect -734 3079 -700 3111
rect -896 3009 -862 3041
rect -896 3007 -862 3009
rect -815 3009 -781 3041
rect -815 3007 -781 3009
rect -734 3009 -700 3041
rect -734 3007 -700 3009
rect -896 2941 -862 2969
rect -896 2935 -862 2941
rect -815 2941 -781 2969
rect -815 2935 -781 2941
rect -734 2941 -700 2969
rect -734 2935 -700 2941
rect -896 2873 -862 2897
rect -896 2863 -862 2873
rect -815 2873 -781 2897
rect -815 2863 -781 2873
rect -734 2873 -700 2897
rect -734 2863 -700 2873
rect -896 2805 -862 2825
rect -896 2791 -862 2805
rect -815 2805 -781 2825
rect -815 2791 -781 2805
rect -734 2805 -700 2825
rect -734 2791 -700 2805
rect -896 2737 -862 2753
rect -896 2719 -862 2737
rect -815 2737 -781 2753
rect -815 2719 -781 2737
rect -734 2737 -700 2753
rect -734 2719 -700 2737
rect -896 2669 -862 2681
rect -896 2647 -862 2669
rect -815 2669 -781 2681
rect -815 2647 -781 2669
rect -734 2669 -700 2681
rect -734 2647 -700 2669
rect -896 2601 -862 2609
rect -896 2575 -862 2601
rect -815 2601 -781 2609
rect -815 2575 -781 2601
rect -734 2601 -700 2609
rect -734 2575 -700 2601
rect -896 2533 -862 2537
rect -896 2503 -862 2533
rect -815 2533 -781 2537
rect -815 2503 -781 2533
rect -734 2533 -700 2537
rect -734 2503 -700 2533
rect -896 2431 -862 2465
rect -815 2431 -781 2465
rect -734 2431 -700 2465
rect -896 2363 -862 2393
rect -896 2359 -862 2363
rect -815 2363 -781 2393
rect -815 2359 -781 2363
rect -734 2363 -700 2393
rect -734 2359 -700 2363
rect -896 2295 -862 2321
rect -896 2287 -862 2295
rect -815 2295 -781 2321
rect -815 2287 -781 2295
rect -734 2295 -700 2321
rect -734 2287 -700 2295
rect -896 2227 -862 2249
rect -896 2215 -862 2227
rect -815 2227 -781 2249
rect -815 2215 -781 2227
rect -734 2227 -700 2249
rect -734 2215 -700 2227
rect -896 2159 -862 2177
rect -896 2143 -862 2159
rect -815 2159 -781 2177
rect -815 2143 -781 2159
rect -734 2159 -700 2177
rect -734 2143 -700 2159
rect -896 2091 -862 2105
rect -896 2071 -862 2091
rect -815 2091 -781 2105
rect -815 2071 -781 2091
rect -734 2091 -700 2105
rect -734 2071 -700 2091
rect -896 2023 -862 2033
rect -896 1999 -862 2023
rect -815 2023 -781 2033
rect -815 1999 -781 2023
rect -734 2023 -700 2033
rect -734 1999 -700 2023
rect -896 1955 -862 1961
rect -896 1927 -862 1955
rect -815 1955 -781 1961
rect -815 1927 -781 1955
rect -734 1955 -700 1961
rect -734 1927 -700 1955
rect -896 1887 -862 1889
rect -896 1855 -862 1887
rect -815 1887 -781 1889
rect -815 1855 -781 1887
rect -734 1887 -700 1889
rect -734 1855 -700 1887
rect -896 1785 -862 1817
rect -896 1783 -862 1785
rect -815 1785 -781 1817
rect -815 1783 -781 1785
rect -734 1785 -700 1817
rect -734 1783 -700 1785
rect -896 1717 -862 1745
rect -896 1711 -862 1717
rect -815 1717 -781 1745
rect -815 1711 -781 1717
rect -734 1717 -700 1745
rect -734 1711 -700 1717
rect -896 1649 -862 1673
rect -896 1639 -862 1649
rect -815 1649 -781 1673
rect -815 1639 -781 1649
rect -734 1649 -700 1673
rect -734 1639 -700 1649
rect -896 1581 -862 1601
rect -896 1567 -862 1581
rect -815 1581 -781 1601
rect -815 1567 -781 1581
rect -734 1581 -700 1601
rect -734 1567 -700 1581
rect -896 1513 -862 1529
rect -896 1495 -862 1513
rect -815 1513 -781 1529
rect -815 1495 -781 1513
rect -734 1513 -700 1529
rect -734 1495 -700 1513
rect -896 1445 -862 1457
rect -896 1423 -862 1445
rect -815 1445 -781 1457
rect -815 1423 -781 1445
rect -734 1445 -700 1457
rect -734 1423 -700 1445
rect -896 1377 -862 1385
rect -896 1351 -862 1377
rect -815 1377 -781 1385
rect -815 1351 -781 1377
rect -734 1377 -700 1385
rect -734 1351 -700 1377
rect -896 1309 -862 1313
rect -896 1279 -862 1309
rect -815 1309 -781 1313
rect -815 1279 -781 1309
rect -734 1309 -700 1313
rect -734 1279 -700 1309
rect -896 1207 -862 1241
rect -815 1207 -781 1241
rect -734 1207 -700 1241
rect -896 1139 -862 1169
rect -896 1135 -862 1139
rect -815 1139 -781 1169
rect -815 1135 -781 1139
rect -734 1139 -700 1169
rect -734 1135 -700 1139
rect -896 1071 -862 1097
rect -896 1063 -862 1071
rect -815 1071 -781 1097
rect -815 1063 -781 1071
rect -734 1071 -700 1097
rect -734 1063 -700 1071
rect -896 1003 -862 1025
rect -896 991 -862 1003
rect -815 1003 -781 1025
rect -815 991 -781 1003
rect -734 1003 -700 1025
rect -734 991 -700 1003
rect -896 935 -862 953
rect -896 919 -862 935
rect -815 935 -781 953
rect -815 919 -781 935
rect -734 935 -700 953
rect -734 919 -700 935
rect -896 867 -862 881
rect -896 847 -862 867
rect -815 867 -781 881
rect -815 847 -781 867
rect -734 867 -700 881
rect -734 847 -700 867
rect -896 799 -862 809
rect -896 775 -862 799
rect -815 799 -781 809
rect -815 775 -781 799
rect -734 799 -700 809
rect -734 775 -700 799
rect -896 731 -862 737
rect -896 703 -862 731
rect -815 731 -781 737
rect -815 703 -781 731
rect -734 731 -700 737
rect -734 703 -700 731
rect -896 663 -862 665
rect -896 631 -862 663
rect -815 663 -781 665
rect -815 631 -781 663
rect -734 663 -700 665
rect -734 631 -700 663
rect -896 561 -862 593
rect -896 559 -862 561
rect -815 561 -781 593
rect -815 559 -781 561
rect -734 561 -700 593
rect -734 559 -700 561
rect -896 493 -862 521
rect -896 487 -862 493
rect -815 493 -781 521
rect -815 487 -781 493
rect -734 493 -700 521
rect -734 487 -700 493
rect -896 425 -862 449
rect -896 415 -862 425
rect -815 425 -781 449
rect -815 415 -781 425
rect -734 425 -700 449
rect -734 415 -700 425
rect -896 357 -862 377
rect -896 343 -862 357
rect -815 357 -781 377
rect -815 343 -781 357
rect -734 357 -700 377
rect -734 343 -700 357
rect -896 289 -862 305
rect -896 271 -862 289
rect -815 289 -781 305
rect -815 271 -781 289
rect -734 289 -700 305
rect -734 271 -700 289
rect -896 221 -862 233
rect -896 199 -862 221
rect -815 221 -781 233
rect -815 199 -781 221
rect -734 221 -700 233
rect -734 199 -700 221
rect -896 153 -862 161
rect -896 127 -862 153
rect -815 153 -781 161
rect -815 127 -781 153
rect -734 153 -700 161
rect -734 127 -700 153
rect -896 85 -862 89
rect -896 55 -862 85
rect -815 85 -781 89
rect -815 55 -781 85
rect -734 85 -700 89
rect -734 55 -700 85
rect -896 -17 -862 17
rect -815 -17 -781 17
rect -734 -17 -700 17
rect -896 -85 -862 -55
rect -896 -89 -862 -85
rect -815 -85 -781 -55
rect -815 -89 -781 -85
rect -734 -85 -700 -55
rect -734 -89 -700 -85
rect -896 -153 -862 -127
rect -896 -161 -862 -153
rect -815 -153 -781 -127
rect -815 -161 -781 -153
rect -734 -153 -700 -127
rect -734 -161 -700 -153
rect -896 -221 -862 -199
rect -896 -233 -862 -221
rect -815 -221 -781 -199
rect -815 -233 -781 -221
rect -734 -221 -700 -199
rect -734 -233 -700 -221
rect -896 -289 -862 -271
rect -896 -305 -862 -289
rect -815 -289 -781 -271
rect -815 -305 -781 -289
rect -734 -289 -700 -271
rect -734 -305 -700 -289
rect -896 -357 -862 -343
rect -896 -377 -862 -357
rect -815 -357 -781 -343
rect -815 -377 -781 -357
rect -734 -357 -700 -343
rect -734 -377 -700 -357
rect -896 -425 -862 -415
rect -896 -449 -862 -425
rect -815 -425 -781 -415
rect -815 -449 -781 -425
rect -734 -425 -700 -415
rect -734 -449 -700 -425
rect -896 -493 -862 -487
rect -896 -521 -862 -493
rect -815 -493 -781 -487
rect -815 -521 -781 -493
rect -734 -493 -700 -487
rect -734 -521 -700 -493
rect -896 -561 -862 -559
rect -896 -593 -862 -561
rect -815 -561 -781 -559
rect -815 -593 -781 -561
rect -734 -561 -700 -559
rect -734 -593 -700 -561
rect -896 -663 -862 -631
rect -896 -665 -862 -663
rect -815 -663 -781 -631
rect -815 -665 -781 -663
rect -734 -663 -700 -631
rect -734 -665 -700 -663
rect -896 -731 -862 -703
rect -896 -737 -862 -731
rect -815 -731 -781 -703
rect -815 -737 -781 -731
rect -734 -731 -700 -703
rect -734 -737 -700 -731
rect -896 -799 -862 -775
rect -896 -809 -862 -799
rect -815 -799 -781 -775
rect -815 -809 -781 -799
rect -734 -799 -700 -775
rect -734 -809 -700 -799
rect -896 -867 -862 -847
rect -896 -881 -862 -867
rect -815 -867 -781 -847
rect -815 -881 -781 -867
rect -734 -867 -700 -847
rect -734 -881 -700 -867
rect -896 -935 -862 -919
rect -896 -953 -862 -935
rect -815 -935 -781 -919
rect -815 -953 -781 -935
rect -734 -935 -700 -919
rect -734 -953 -700 -935
rect -896 -1003 -862 -991
rect -896 -1025 -862 -1003
rect -815 -1003 -781 -991
rect -815 -1025 -781 -1003
rect -734 -1003 -700 -991
rect -734 -1025 -700 -1003
rect -896 -1071 -862 -1063
rect -896 -1097 -862 -1071
rect -815 -1071 -781 -1063
rect -815 -1097 -781 -1071
rect -734 -1071 -700 -1063
rect -734 -1097 -700 -1071
rect -896 -1139 -862 -1135
rect -896 -1169 -862 -1139
rect -815 -1139 -781 -1135
rect -815 -1169 -781 -1139
rect -734 -1139 -700 -1135
rect -734 -1169 -700 -1139
rect -896 -1241 -862 -1207
rect -815 -1241 -781 -1207
rect -734 -1241 -700 -1207
rect -896 -1309 -862 -1279
rect -896 -1313 -862 -1309
rect -815 -1309 -781 -1279
rect -815 -1313 -781 -1309
rect -734 -1309 -700 -1279
rect -734 -1313 -700 -1309
rect -896 -1377 -862 -1351
rect -896 -1385 -862 -1377
rect -815 -1377 -781 -1351
rect -815 -1385 -781 -1377
rect -734 -1377 -700 -1351
rect -734 -1385 -700 -1377
rect -896 -1445 -862 -1423
rect -896 -1457 -862 -1445
rect -815 -1445 -781 -1423
rect -815 -1457 -781 -1445
rect -734 -1445 -700 -1423
rect -734 -1457 -700 -1445
rect -896 -1513 -862 -1495
rect -896 -1529 -862 -1513
rect -815 -1513 -781 -1495
rect -815 -1529 -781 -1513
rect -734 -1513 -700 -1495
rect -734 -1529 -700 -1513
rect -896 -1581 -862 -1567
rect -896 -1601 -862 -1581
rect -815 -1581 -781 -1567
rect -815 -1601 -781 -1581
rect -734 -1581 -700 -1567
rect -734 -1601 -700 -1581
rect -896 -1649 -862 -1639
rect -896 -1673 -862 -1649
rect -815 -1649 -781 -1639
rect -815 -1673 -781 -1649
rect -734 -1649 -700 -1639
rect -734 -1673 -700 -1649
rect -896 -1717 -862 -1711
rect -896 -1745 -862 -1717
rect -815 -1717 -781 -1711
rect -815 -1745 -781 -1717
rect -734 -1717 -700 -1711
rect -734 -1745 -700 -1717
rect -896 -1785 -862 -1783
rect -896 -1817 -862 -1785
rect -815 -1785 -781 -1783
rect -815 -1817 -781 -1785
rect -734 -1785 -700 -1783
rect -734 -1817 -700 -1785
rect -896 -1887 -862 -1855
rect -896 -1889 -862 -1887
rect -815 -1887 -781 -1855
rect -815 -1889 -781 -1887
rect -734 -1887 -700 -1855
rect -734 -1889 -700 -1887
rect -896 -1955 -862 -1927
rect -896 -1961 -862 -1955
rect -815 -1955 -781 -1927
rect -815 -1961 -781 -1955
rect -734 -1955 -700 -1927
rect -734 -1961 -700 -1955
rect -896 -2023 -862 -1999
rect -896 -2033 -862 -2023
rect -815 -2023 -781 -1999
rect -815 -2033 -781 -2023
rect -734 -2023 -700 -1999
rect -734 -2033 -700 -2023
rect -896 -2091 -862 -2071
rect -896 -2105 -862 -2091
rect -815 -2091 -781 -2071
rect -815 -2105 -781 -2091
rect -734 -2091 -700 -2071
rect -734 -2105 -700 -2091
rect -896 -2159 -862 -2143
rect -896 -2177 -862 -2159
rect -815 -2159 -781 -2143
rect -815 -2177 -781 -2159
rect -734 -2159 -700 -2143
rect -734 -2177 -700 -2159
rect -896 -2227 -862 -2215
rect -896 -2249 -862 -2227
rect -815 -2227 -781 -2215
rect -815 -2249 -781 -2227
rect -734 -2227 -700 -2215
rect -734 -2249 -700 -2227
rect -896 -2295 -862 -2287
rect -896 -2321 -862 -2295
rect -815 -2295 -781 -2287
rect -815 -2321 -781 -2295
rect -734 -2295 -700 -2287
rect -734 -2321 -700 -2295
rect -896 -2363 -862 -2359
rect -896 -2393 -862 -2363
rect -815 -2363 -781 -2359
rect -815 -2393 -781 -2363
rect -734 -2363 -700 -2359
rect -734 -2393 -700 -2363
rect -896 -2465 -862 -2431
rect -815 -2465 -781 -2431
rect -734 -2465 -700 -2431
rect -896 -2533 -862 -2503
rect -896 -2537 -862 -2533
rect -815 -2533 -781 -2503
rect -815 -2537 -781 -2533
rect -734 -2533 -700 -2503
rect -734 -2537 -700 -2533
rect -896 -2601 -862 -2575
rect -896 -2609 -862 -2601
rect -815 -2601 -781 -2575
rect -815 -2609 -781 -2601
rect -734 -2601 -700 -2575
rect -734 -2609 -700 -2601
rect -896 -2669 -862 -2647
rect -896 -2681 -862 -2669
rect -815 -2669 -781 -2647
rect -815 -2681 -781 -2669
rect -734 -2669 -700 -2647
rect -734 -2681 -700 -2669
rect -896 -2737 -862 -2719
rect -896 -2753 -862 -2737
rect -815 -2737 -781 -2719
rect -815 -2753 -781 -2737
rect -734 -2737 -700 -2719
rect -734 -2753 -700 -2737
rect -896 -2805 -862 -2791
rect -896 -2825 -862 -2805
rect -815 -2805 -781 -2791
rect -815 -2825 -781 -2805
rect -734 -2805 -700 -2791
rect -734 -2825 -700 -2805
rect -896 -2873 -862 -2863
rect -896 -2897 -862 -2873
rect -815 -2873 -781 -2863
rect -815 -2897 -781 -2873
rect -734 -2873 -700 -2863
rect -734 -2897 -700 -2873
rect -896 -2941 -862 -2935
rect -896 -2969 -862 -2941
rect -815 -2941 -781 -2935
rect -815 -2969 -781 -2941
rect -734 -2941 -700 -2935
rect -734 -2969 -700 -2941
rect -896 -3009 -862 -3007
rect -896 -3041 -862 -3009
rect -815 -3009 -781 -3007
rect -815 -3041 -781 -3009
rect -734 -3009 -700 -3007
rect -734 -3041 -700 -3009
rect -896 -3111 -862 -3079
rect -896 -3113 -862 -3111
rect -815 -3111 -781 -3079
rect -815 -3113 -781 -3111
rect -734 -3111 -700 -3079
rect -734 -3113 -700 -3111
rect -896 -3179 -862 -3151
rect -896 -3185 -862 -3179
rect -815 -3179 -781 -3151
rect -815 -3185 -781 -3179
rect -734 -3179 -700 -3151
rect -734 -3185 -700 -3179
rect -896 -3247 -862 -3223
rect -896 -3257 -862 -3247
rect -815 -3247 -781 -3223
rect -815 -3257 -781 -3247
rect -734 -3247 -700 -3223
rect -734 -3257 -700 -3247
rect -896 -3315 -862 -3295
rect -896 -3329 -862 -3315
rect -815 -3315 -781 -3295
rect -815 -3329 -781 -3315
rect -734 -3315 -700 -3295
rect -734 -3329 -700 -3315
rect -896 -3383 -862 -3367
rect -896 -3401 -862 -3383
rect -815 -3383 -781 -3367
rect -815 -3401 -781 -3383
rect -734 -3383 -700 -3367
rect -734 -3401 -700 -3383
rect -896 -3451 -862 -3439
rect -896 -3473 -862 -3451
rect -815 -3451 -781 -3439
rect -815 -3473 -781 -3451
rect -734 -3451 -700 -3439
rect -734 -3473 -700 -3451
rect -896 -3519 -862 -3511
rect -896 -3545 -862 -3519
rect -815 -3519 -781 -3511
rect -815 -3545 -781 -3519
rect -734 -3519 -700 -3511
rect -734 -3545 -700 -3519
rect -896 -3587 -862 -3583
rect -896 -3617 -862 -3587
rect -815 -3587 -781 -3583
rect -815 -3617 -781 -3587
rect -734 -3587 -700 -3583
rect -734 -3617 -700 -3587
rect -896 -3689 -862 -3655
rect -815 -3689 -781 -3655
rect -734 -3689 -700 -3655
rect -896 -3757 -862 -3727
rect -896 -3761 -862 -3757
rect -815 -3757 -781 -3727
rect -815 -3761 -781 -3757
rect -734 -3757 -700 -3727
rect -734 -3761 -700 -3757
rect -896 -3825 -862 -3799
rect -896 -3833 -862 -3825
rect -815 -3825 -781 -3799
rect -815 -3833 -781 -3825
rect -734 -3825 -700 -3799
rect -734 -3833 -700 -3825
rect -896 -3893 -862 -3871
rect -896 -3905 -862 -3893
rect -815 -3893 -781 -3871
rect -815 -3905 -781 -3893
rect -734 -3893 -700 -3871
rect -734 -3905 -700 -3893
rect -896 -3961 -862 -3943
rect -896 -3977 -862 -3961
rect -815 -3961 -781 -3943
rect -815 -3977 -781 -3961
rect -734 -3961 -700 -3943
rect -734 -3977 -700 -3961
rect -896 -4029 -862 -4015
rect -896 -4049 -862 -4029
rect -815 -4029 -781 -4015
rect -815 -4049 -781 -4029
rect -734 -4029 -700 -4015
rect -734 -4049 -700 -4029
rect -896 -4097 -862 -4087
rect -896 -4121 -862 -4097
rect -815 -4097 -781 -4087
rect -815 -4121 -781 -4097
rect -734 -4097 -700 -4087
rect -734 -4121 -700 -4097
rect -896 -4165 -862 -4159
rect -896 -4193 -862 -4165
rect -815 -4165 -781 -4159
rect -815 -4193 -781 -4165
rect -734 -4165 -700 -4159
rect -734 -4193 -700 -4165
rect -896 -4233 -862 -4231
rect -896 -4265 -862 -4233
rect -815 -4233 -781 -4231
rect -815 -4265 -781 -4233
rect -734 -4233 -700 -4231
rect -734 -4265 -700 -4233
rect -896 -4335 -862 -4303
rect -896 -4337 -862 -4335
rect -815 -4335 -781 -4303
rect -815 -4337 -781 -4335
rect -734 -4335 -700 -4303
rect -734 -4337 -700 -4335
rect -896 -4403 -862 -4375
rect -896 -4409 -862 -4403
rect -815 -4403 -781 -4375
rect -815 -4409 -781 -4403
rect -734 -4403 -700 -4375
rect -734 -4409 -700 -4403
rect -896 -4471 -862 -4447
rect -896 -4481 -862 -4471
rect -815 -4471 -781 -4447
rect -815 -4481 -781 -4471
rect -734 -4471 -700 -4447
rect -734 -4481 -700 -4471
rect -896 -4539 -862 -4519
rect -896 -4553 -862 -4539
rect -815 -4539 -781 -4519
rect -815 -4553 -781 -4539
rect -734 -4539 -700 -4519
rect -734 -4553 -700 -4539
rect -896 -4607 -862 -4591
rect -896 -4625 -862 -4607
rect -815 -4607 -781 -4591
rect -815 -4625 -781 -4607
rect -734 -4607 -700 -4591
rect -734 -4625 -700 -4607
rect -896 -4675 -862 -4663
rect -896 -4697 -862 -4675
rect -815 -4675 -781 -4663
rect -815 -4697 -781 -4675
rect -734 -4675 -700 -4663
rect -734 -4697 -700 -4675
rect -896 -4743 -862 -4735
rect -896 -4769 -862 -4743
rect -815 -4743 -781 -4735
rect -815 -4769 -781 -4743
rect -734 -4743 -700 -4735
rect -734 -4769 -700 -4743
rect -896 -4811 -862 -4807
rect -896 -4841 -862 -4811
rect -815 -4811 -781 -4807
rect -815 -4841 -781 -4811
rect -734 -4811 -700 -4807
rect -734 -4841 -700 -4811
rect -896 -4913 -862 -4879
rect -815 -4913 -781 -4879
rect -734 -4913 -700 -4879
rect -896 -4981 -862 -4951
rect -896 -4985 -862 -4981
rect -815 -4981 -781 -4951
rect -815 -4985 -781 -4981
rect -734 -4981 -700 -4951
rect -734 -4985 -700 -4981
rect -585 4981 -479 4985
rect -585 -4981 -479 4981
rect -585 -4985 -479 -4981
rect -364 4981 -330 4985
rect -364 4951 -330 4981
rect -283 4981 -249 4985
rect -283 4951 -249 4981
rect -202 4981 -168 4985
rect -202 4951 -168 4981
rect -364 4879 -330 4913
rect -283 4879 -249 4913
rect -202 4879 -168 4913
rect -364 4811 -330 4841
rect -364 4807 -330 4811
rect -283 4811 -249 4841
rect -283 4807 -249 4811
rect -202 4811 -168 4841
rect -202 4807 -168 4811
rect -364 4743 -330 4769
rect -364 4735 -330 4743
rect -283 4743 -249 4769
rect -283 4735 -249 4743
rect -202 4743 -168 4769
rect -202 4735 -168 4743
rect -364 4675 -330 4697
rect -364 4663 -330 4675
rect -283 4675 -249 4697
rect -283 4663 -249 4675
rect -202 4675 -168 4697
rect -202 4663 -168 4675
rect -364 4607 -330 4625
rect -364 4591 -330 4607
rect -283 4607 -249 4625
rect -283 4591 -249 4607
rect -202 4607 -168 4625
rect -202 4591 -168 4607
rect -364 4539 -330 4553
rect -364 4519 -330 4539
rect -283 4539 -249 4553
rect -283 4519 -249 4539
rect -202 4539 -168 4553
rect -202 4519 -168 4539
rect -364 4471 -330 4481
rect -364 4447 -330 4471
rect -283 4471 -249 4481
rect -283 4447 -249 4471
rect -202 4471 -168 4481
rect -202 4447 -168 4471
rect -364 4403 -330 4409
rect -364 4375 -330 4403
rect -283 4403 -249 4409
rect -283 4375 -249 4403
rect -202 4403 -168 4409
rect -202 4375 -168 4403
rect -364 4335 -330 4337
rect -364 4303 -330 4335
rect -283 4335 -249 4337
rect -283 4303 -249 4335
rect -202 4335 -168 4337
rect -202 4303 -168 4335
rect -364 4233 -330 4265
rect -364 4231 -330 4233
rect -283 4233 -249 4265
rect -283 4231 -249 4233
rect -202 4233 -168 4265
rect -202 4231 -168 4233
rect -364 4165 -330 4193
rect -364 4159 -330 4165
rect -283 4165 -249 4193
rect -283 4159 -249 4165
rect -202 4165 -168 4193
rect -202 4159 -168 4165
rect -364 4097 -330 4121
rect -364 4087 -330 4097
rect -283 4097 -249 4121
rect -283 4087 -249 4097
rect -202 4097 -168 4121
rect -202 4087 -168 4097
rect -364 4029 -330 4049
rect -364 4015 -330 4029
rect -283 4029 -249 4049
rect -283 4015 -249 4029
rect -202 4029 -168 4049
rect -202 4015 -168 4029
rect -364 3961 -330 3977
rect -364 3943 -330 3961
rect -283 3961 -249 3977
rect -283 3943 -249 3961
rect -202 3961 -168 3977
rect -202 3943 -168 3961
rect -364 3893 -330 3905
rect -364 3871 -330 3893
rect -283 3893 -249 3905
rect -283 3871 -249 3893
rect -202 3893 -168 3905
rect -202 3871 -168 3893
rect -364 3825 -330 3833
rect -364 3799 -330 3825
rect -283 3825 -249 3833
rect -283 3799 -249 3825
rect -202 3825 -168 3833
rect -202 3799 -168 3825
rect -364 3757 -330 3761
rect -364 3727 -330 3757
rect -283 3757 -249 3761
rect -283 3727 -249 3757
rect -202 3757 -168 3761
rect -202 3727 -168 3757
rect -364 3655 -330 3689
rect -283 3655 -249 3689
rect -202 3655 -168 3689
rect -364 3587 -330 3617
rect -364 3583 -330 3587
rect -283 3587 -249 3617
rect -283 3583 -249 3587
rect -202 3587 -168 3617
rect -202 3583 -168 3587
rect -364 3519 -330 3545
rect -364 3511 -330 3519
rect -283 3519 -249 3545
rect -283 3511 -249 3519
rect -202 3519 -168 3545
rect -202 3511 -168 3519
rect -364 3451 -330 3473
rect -364 3439 -330 3451
rect -283 3451 -249 3473
rect -283 3439 -249 3451
rect -202 3451 -168 3473
rect -202 3439 -168 3451
rect -364 3383 -330 3401
rect -364 3367 -330 3383
rect -283 3383 -249 3401
rect -283 3367 -249 3383
rect -202 3383 -168 3401
rect -202 3367 -168 3383
rect -364 3315 -330 3329
rect -364 3295 -330 3315
rect -283 3315 -249 3329
rect -283 3295 -249 3315
rect -202 3315 -168 3329
rect -202 3295 -168 3315
rect -364 3247 -330 3257
rect -364 3223 -330 3247
rect -283 3247 -249 3257
rect -283 3223 -249 3247
rect -202 3247 -168 3257
rect -202 3223 -168 3247
rect -364 3179 -330 3185
rect -364 3151 -330 3179
rect -283 3179 -249 3185
rect -283 3151 -249 3179
rect -202 3179 -168 3185
rect -202 3151 -168 3179
rect -364 3111 -330 3113
rect -364 3079 -330 3111
rect -283 3111 -249 3113
rect -283 3079 -249 3111
rect -202 3111 -168 3113
rect -202 3079 -168 3111
rect -364 3009 -330 3041
rect -364 3007 -330 3009
rect -283 3009 -249 3041
rect -283 3007 -249 3009
rect -202 3009 -168 3041
rect -202 3007 -168 3009
rect -364 2941 -330 2969
rect -364 2935 -330 2941
rect -283 2941 -249 2969
rect -283 2935 -249 2941
rect -202 2941 -168 2969
rect -202 2935 -168 2941
rect -364 2873 -330 2897
rect -364 2863 -330 2873
rect -283 2873 -249 2897
rect -283 2863 -249 2873
rect -202 2873 -168 2897
rect -202 2863 -168 2873
rect -364 2805 -330 2825
rect -364 2791 -330 2805
rect -283 2805 -249 2825
rect -283 2791 -249 2805
rect -202 2805 -168 2825
rect -202 2791 -168 2805
rect -364 2737 -330 2753
rect -364 2719 -330 2737
rect -283 2737 -249 2753
rect -283 2719 -249 2737
rect -202 2737 -168 2753
rect -202 2719 -168 2737
rect -364 2669 -330 2681
rect -364 2647 -330 2669
rect -283 2669 -249 2681
rect -283 2647 -249 2669
rect -202 2669 -168 2681
rect -202 2647 -168 2669
rect -364 2601 -330 2609
rect -364 2575 -330 2601
rect -283 2601 -249 2609
rect -283 2575 -249 2601
rect -202 2601 -168 2609
rect -202 2575 -168 2601
rect -364 2533 -330 2537
rect -364 2503 -330 2533
rect -283 2533 -249 2537
rect -283 2503 -249 2533
rect -202 2533 -168 2537
rect -202 2503 -168 2533
rect -364 2431 -330 2465
rect -283 2431 -249 2465
rect -202 2431 -168 2465
rect -364 2363 -330 2393
rect -364 2359 -330 2363
rect -283 2363 -249 2393
rect -283 2359 -249 2363
rect -202 2363 -168 2393
rect -202 2359 -168 2363
rect -364 2295 -330 2321
rect -364 2287 -330 2295
rect -283 2295 -249 2321
rect -283 2287 -249 2295
rect -202 2295 -168 2321
rect -202 2287 -168 2295
rect -364 2227 -330 2249
rect -364 2215 -330 2227
rect -283 2227 -249 2249
rect -283 2215 -249 2227
rect -202 2227 -168 2249
rect -202 2215 -168 2227
rect -364 2159 -330 2177
rect -364 2143 -330 2159
rect -283 2159 -249 2177
rect -283 2143 -249 2159
rect -202 2159 -168 2177
rect -202 2143 -168 2159
rect -364 2091 -330 2105
rect -364 2071 -330 2091
rect -283 2091 -249 2105
rect -283 2071 -249 2091
rect -202 2091 -168 2105
rect -202 2071 -168 2091
rect -364 2023 -330 2033
rect -364 1999 -330 2023
rect -283 2023 -249 2033
rect -283 1999 -249 2023
rect -202 2023 -168 2033
rect -202 1999 -168 2023
rect -364 1955 -330 1961
rect -364 1927 -330 1955
rect -283 1955 -249 1961
rect -283 1927 -249 1955
rect -202 1955 -168 1961
rect -202 1927 -168 1955
rect -364 1887 -330 1889
rect -364 1855 -330 1887
rect -283 1887 -249 1889
rect -283 1855 -249 1887
rect -202 1887 -168 1889
rect -202 1855 -168 1887
rect -364 1785 -330 1817
rect -364 1783 -330 1785
rect -283 1785 -249 1817
rect -283 1783 -249 1785
rect -202 1785 -168 1817
rect -202 1783 -168 1785
rect -364 1717 -330 1745
rect -364 1711 -330 1717
rect -283 1717 -249 1745
rect -283 1711 -249 1717
rect -202 1717 -168 1745
rect -202 1711 -168 1717
rect -364 1649 -330 1673
rect -364 1639 -330 1649
rect -283 1649 -249 1673
rect -283 1639 -249 1649
rect -202 1649 -168 1673
rect -202 1639 -168 1649
rect -364 1581 -330 1601
rect -364 1567 -330 1581
rect -283 1581 -249 1601
rect -283 1567 -249 1581
rect -202 1581 -168 1601
rect -202 1567 -168 1581
rect -364 1513 -330 1529
rect -364 1495 -330 1513
rect -283 1513 -249 1529
rect -283 1495 -249 1513
rect -202 1513 -168 1529
rect -202 1495 -168 1513
rect -364 1445 -330 1457
rect -364 1423 -330 1445
rect -283 1445 -249 1457
rect -283 1423 -249 1445
rect -202 1445 -168 1457
rect -202 1423 -168 1445
rect -364 1377 -330 1385
rect -364 1351 -330 1377
rect -283 1377 -249 1385
rect -283 1351 -249 1377
rect -202 1377 -168 1385
rect -202 1351 -168 1377
rect -364 1309 -330 1313
rect -364 1279 -330 1309
rect -283 1309 -249 1313
rect -283 1279 -249 1309
rect -202 1309 -168 1313
rect -202 1279 -168 1309
rect -364 1207 -330 1241
rect -283 1207 -249 1241
rect -202 1207 -168 1241
rect -364 1139 -330 1169
rect -364 1135 -330 1139
rect -283 1139 -249 1169
rect -283 1135 -249 1139
rect -202 1139 -168 1169
rect -202 1135 -168 1139
rect -364 1071 -330 1097
rect -364 1063 -330 1071
rect -283 1071 -249 1097
rect -283 1063 -249 1071
rect -202 1071 -168 1097
rect -202 1063 -168 1071
rect -364 1003 -330 1025
rect -364 991 -330 1003
rect -283 1003 -249 1025
rect -283 991 -249 1003
rect -202 1003 -168 1025
rect -202 991 -168 1003
rect -364 935 -330 953
rect -364 919 -330 935
rect -283 935 -249 953
rect -283 919 -249 935
rect -202 935 -168 953
rect -202 919 -168 935
rect -364 867 -330 881
rect -364 847 -330 867
rect -283 867 -249 881
rect -283 847 -249 867
rect -202 867 -168 881
rect -202 847 -168 867
rect -364 799 -330 809
rect -364 775 -330 799
rect -283 799 -249 809
rect -283 775 -249 799
rect -202 799 -168 809
rect -202 775 -168 799
rect -364 731 -330 737
rect -364 703 -330 731
rect -283 731 -249 737
rect -283 703 -249 731
rect -202 731 -168 737
rect -202 703 -168 731
rect -364 663 -330 665
rect -364 631 -330 663
rect -283 663 -249 665
rect -283 631 -249 663
rect -202 663 -168 665
rect -202 631 -168 663
rect -364 561 -330 593
rect -364 559 -330 561
rect -283 561 -249 593
rect -283 559 -249 561
rect -202 561 -168 593
rect -202 559 -168 561
rect -364 493 -330 521
rect -364 487 -330 493
rect -283 493 -249 521
rect -283 487 -249 493
rect -202 493 -168 521
rect -202 487 -168 493
rect -364 425 -330 449
rect -364 415 -330 425
rect -283 425 -249 449
rect -283 415 -249 425
rect -202 425 -168 449
rect -202 415 -168 425
rect -364 357 -330 377
rect -364 343 -330 357
rect -283 357 -249 377
rect -283 343 -249 357
rect -202 357 -168 377
rect -202 343 -168 357
rect -364 289 -330 305
rect -364 271 -330 289
rect -283 289 -249 305
rect -283 271 -249 289
rect -202 289 -168 305
rect -202 271 -168 289
rect -364 221 -330 233
rect -364 199 -330 221
rect -283 221 -249 233
rect -283 199 -249 221
rect -202 221 -168 233
rect -202 199 -168 221
rect -364 153 -330 161
rect -364 127 -330 153
rect -283 153 -249 161
rect -283 127 -249 153
rect -202 153 -168 161
rect -202 127 -168 153
rect -364 85 -330 89
rect -364 55 -330 85
rect -283 85 -249 89
rect -283 55 -249 85
rect -202 85 -168 89
rect -202 55 -168 85
rect -364 -17 -330 17
rect -283 -17 -249 17
rect -202 -17 -168 17
rect -364 -85 -330 -55
rect -364 -89 -330 -85
rect -283 -85 -249 -55
rect -283 -89 -249 -85
rect -202 -85 -168 -55
rect -202 -89 -168 -85
rect -364 -153 -330 -127
rect -364 -161 -330 -153
rect -283 -153 -249 -127
rect -283 -161 -249 -153
rect -202 -153 -168 -127
rect -202 -161 -168 -153
rect -364 -221 -330 -199
rect -364 -233 -330 -221
rect -283 -221 -249 -199
rect -283 -233 -249 -221
rect -202 -221 -168 -199
rect -202 -233 -168 -221
rect -364 -289 -330 -271
rect -364 -305 -330 -289
rect -283 -289 -249 -271
rect -283 -305 -249 -289
rect -202 -289 -168 -271
rect -202 -305 -168 -289
rect -364 -357 -330 -343
rect -364 -377 -330 -357
rect -283 -357 -249 -343
rect -283 -377 -249 -357
rect -202 -357 -168 -343
rect -202 -377 -168 -357
rect -364 -425 -330 -415
rect -364 -449 -330 -425
rect -283 -425 -249 -415
rect -283 -449 -249 -425
rect -202 -425 -168 -415
rect -202 -449 -168 -425
rect -364 -493 -330 -487
rect -364 -521 -330 -493
rect -283 -493 -249 -487
rect -283 -521 -249 -493
rect -202 -493 -168 -487
rect -202 -521 -168 -493
rect -364 -561 -330 -559
rect -364 -593 -330 -561
rect -283 -561 -249 -559
rect -283 -593 -249 -561
rect -202 -561 -168 -559
rect -202 -593 -168 -561
rect -364 -663 -330 -631
rect -364 -665 -330 -663
rect -283 -663 -249 -631
rect -283 -665 -249 -663
rect -202 -663 -168 -631
rect -202 -665 -168 -663
rect -364 -731 -330 -703
rect -364 -737 -330 -731
rect -283 -731 -249 -703
rect -283 -737 -249 -731
rect -202 -731 -168 -703
rect -202 -737 -168 -731
rect -364 -799 -330 -775
rect -364 -809 -330 -799
rect -283 -799 -249 -775
rect -283 -809 -249 -799
rect -202 -799 -168 -775
rect -202 -809 -168 -799
rect -364 -867 -330 -847
rect -364 -881 -330 -867
rect -283 -867 -249 -847
rect -283 -881 -249 -867
rect -202 -867 -168 -847
rect -202 -881 -168 -867
rect -364 -935 -330 -919
rect -364 -953 -330 -935
rect -283 -935 -249 -919
rect -283 -953 -249 -935
rect -202 -935 -168 -919
rect -202 -953 -168 -935
rect -364 -1003 -330 -991
rect -364 -1025 -330 -1003
rect -283 -1003 -249 -991
rect -283 -1025 -249 -1003
rect -202 -1003 -168 -991
rect -202 -1025 -168 -1003
rect -364 -1071 -330 -1063
rect -364 -1097 -330 -1071
rect -283 -1071 -249 -1063
rect -283 -1097 -249 -1071
rect -202 -1071 -168 -1063
rect -202 -1097 -168 -1071
rect -364 -1139 -330 -1135
rect -364 -1169 -330 -1139
rect -283 -1139 -249 -1135
rect -283 -1169 -249 -1139
rect -202 -1139 -168 -1135
rect -202 -1169 -168 -1139
rect -364 -1241 -330 -1207
rect -283 -1241 -249 -1207
rect -202 -1241 -168 -1207
rect -364 -1309 -330 -1279
rect -364 -1313 -330 -1309
rect -283 -1309 -249 -1279
rect -283 -1313 -249 -1309
rect -202 -1309 -168 -1279
rect -202 -1313 -168 -1309
rect -364 -1377 -330 -1351
rect -364 -1385 -330 -1377
rect -283 -1377 -249 -1351
rect -283 -1385 -249 -1377
rect -202 -1377 -168 -1351
rect -202 -1385 -168 -1377
rect -364 -1445 -330 -1423
rect -364 -1457 -330 -1445
rect -283 -1445 -249 -1423
rect -283 -1457 -249 -1445
rect -202 -1445 -168 -1423
rect -202 -1457 -168 -1445
rect -364 -1513 -330 -1495
rect -364 -1529 -330 -1513
rect -283 -1513 -249 -1495
rect -283 -1529 -249 -1513
rect -202 -1513 -168 -1495
rect -202 -1529 -168 -1513
rect -364 -1581 -330 -1567
rect -364 -1601 -330 -1581
rect -283 -1581 -249 -1567
rect -283 -1601 -249 -1581
rect -202 -1581 -168 -1567
rect -202 -1601 -168 -1581
rect -364 -1649 -330 -1639
rect -364 -1673 -330 -1649
rect -283 -1649 -249 -1639
rect -283 -1673 -249 -1649
rect -202 -1649 -168 -1639
rect -202 -1673 -168 -1649
rect -364 -1717 -330 -1711
rect -364 -1745 -330 -1717
rect -283 -1717 -249 -1711
rect -283 -1745 -249 -1717
rect -202 -1717 -168 -1711
rect -202 -1745 -168 -1717
rect -364 -1785 -330 -1783
rect -364 -1817 -330 -1785
rect -283 -1785 -249 -1783
rect -283 -1817 -249 -1785
rect -202 -1785 -168 -1783
rect -202 -1817 -168 -1785
rect -364 -1887 -330 -1855
rect -364 -1889 -330 -1887
rect -283 -1887 -249 -1855
rect -283 -1889 -249 -1887
rect -202 -1887 -168 -1855
rect -202 -1889 -168 -1887
rect -364 -1955 -330 -1927
rect -364 -1961 -330 -1955
rect -283 -1955 -249 -1927
rect -283 -1961 -249 -1955
rect -202 -1955 -168 -1927
rect -202 -1961 -168 -1955
rect -364 -2023 -330 -1999
rect -364 -2033 -330 -2023
rect -283 -2023 -249 -1999
rect -283 -2033 -249 -2023
rect -202 -2023 -168 -1999
rect -202 -2033 -168 -2023
rect -364 -2091 -330 -2071
rect -364 -2105 -330 -2091
rect -283 -2091 -249 -2071
rect -283 -2105 -249 -2091
rect -202 -2091 -168 -2071
rect -202 -2105 -168 -2091
rect -364 -2159 -330 -2143
rect -364 -2177 -330 -2159
rect -283 -2159 -249 -2143
rect -283 -2177 -249 -2159
rect -202 -2159 -168 -2143
rect -202 -2177 -168 -2159
rect -364 -2227 -330 -2215
rect -364 -2249 -330 -2227
rect -283 -2227 -249 -2215
rect -283 -2249 -249 -2227
rect -202 -2227 -168 -2215
rect -202 -2249 -168 -2227
rect -364 -2295 -330 -2287
rect -364 -2321 -330 -2295
rect -283 -2295 -249 -2287
rect -283 -2321 -249 -2295
rect -202 -2295 -168 -2287
rect -202 -2321 -168 -2295
rect -364 -2363 -330 -2359
rect -364 -2393 -330 -2363
rect -283 -2363 -249 -2359
rect -283 -2393 -249 -2363
rect -202 -2363 -168 -2359
rect -202 -2393 -168 -2363
rect -364 -2465 -330 -2431
rect -283 -2465 -249 -2431
rect -202 -2465 -168 -2431
rect -364 -2533 -330 -2503
rect -364 -2537 -330 -2533
rect -283 -2533 -249 -2503
rect -283 -2537 -249 -2533
rect -202 -2533 -168 -2503
rect -202 -2537 -168 -2533
rect -364 -2601 -330 -2575
rect -364 -2609 -330 -2601
rect -283 -2601 -249 -2575
rect -283 -2609 -249 -2601
rect -202 -2601 -168 -2575
rect -202 -2609 -168 -2601
rect -364 -2669 -330 -2647
rect -364 -2681 -330 -2669
rect -283 -2669 -249 -2647
rect -283 -2681 -249 -2669
rect -202 -2669 -168 -2647
rect -202 -2681 -168 -2669
rect -364 -2737 -330 -2719
rect -364 -2753 -330 -2737
rect -283 -2737 -249 -2719
rect -283 -2753 -249 -2737
rect -202 -2737 -168 -2719
rect -202 -2753 -168 -2737
rect -364 -2805 -330 -2791
rect -364 -2825 -330 -2805
rect -283 -2805 -249 -2791
rect -283 -2825 -249 -2805
rect -202 -2805 -168 -2791
rect -202 -2825 -168 -2805
rect -364 -2873 -330 -2863
rect -364 -2897 -330 -2873
rect -283 -2873 -249 -2863
rect -283 -2897 -249 -2873
rect -202 -2873 -168 -2863
rect -202 -2897 -168 -2873
rect -364 -2941 -330 -2935
rect -364 -2969 -330 -2941
rect -283 -2941 -249 -2935
rect -283 -2969 -249 -2941
rect -202 -2941 -168 -2935
rect -202 -2969 -168 -2941
rect -364 -3009 -330 -3007
rect -364 -3041 -330 -3009
rect -283 -3009 -249 -3007
rect -283 -3041 -249 -3009
rect -202 -3009 -168 -3007
rect -202 -3041 -168 -3009
rect -364 -3111 -330 -3079
rect -364 -3113 -330 -3111
rect -283 -3111 -249 -3079
rect -283 -3113 -249 -3111
rect -202 -3111 -168 -3079
rect -202 -3113 -168 -3111
rect -364 -3179 -330 -3151
rect -364 -3185 -330 -3179
rect -283 -3179 -249 -3151
rect -283 -3185 -249 -3179
rect -202 -3179 -168 -3151
rect -202 -3185 -168 -3179
rect -364 -3247 -330 -3223
rect -364 -3257 -330 -3247
rect -283 -3247 -249 -3223
rect -283 -3257 -249 -3247
rect -202 -3247 -168 -3223
rect -202 -3257 -168 -3247
rect -364 -3315 -330 -3295
rect -364 -3329 -330 -3315
rect -283 -3315 -249 -3295
rect -283 -3329 -249 -3315
rect -202 -3315 -168 -3295
rect -202 -3329 -168 -3315
rect -364 -3383 -330 -3367
rect -364 -3401 -330 -3383
rect -283 -3383 -249 -3367
rect -283 -3401 -249 -3383
rect -202 -3383 -168 -3367
rect -202 -3401 -168 -3383
rect -364 -3451 -330 -3439
rect -364 -3473 -330 -3451
rect -283 -3451 -249 -3439
rect -283 -3473 -249 -3451
rect -202 -3451 -168 -3439
rect -202 -3473 -168 -3451
rect -364 -3519 -330 -3511
rect -364 -3545 -330 -3519
rect -283 -3519 -249 -3511
rect -283 -3545 -249 -3519
rect -202 -3519 -168 -3511
rect -202 -3545 -168 -3519
rect -364 -3587 -330 -3583
rect -364 -3617 -330 -3587
rect -283 -3587 -249 -3583
rect -283 -3617 -249 -3587
rect -202 -3587 -168 -3583
rect -202 -3617 -168 -3587
rect -364 -3689 -330 -3655
rect -283 -3689 -249 -3655
rect -202 -3689 -168 -3655
rect -364 -3757 -330 -3727
rect -364 -3761 -330 -3757
rect -283 -3757 -249 -3727
rect -283 -3761 -249 -3757
rect -202 -3757 -168 -3727
rect -202 -3761 -168 -3757
rect -364 -3825 -330 -3799
rect -364 -3833 -330 -3825
rect -283 -3825 -249 -3799
rect -283 -3833 -249 -3825
rect -202 -3825 -168 -3799
rect -202 -3833 -168 -3825
rect -364 -3893 -330 -3871
rect -364 -3905 -330 -3893
rect -283 -3893 -249 -3871
rect -283 -3905 -249 -3893
rect -202 -3893 -168 -3871
rect -202 -3905 -168 -3893
rect -364 -3961 -330 -3943
rect -364 -3977 -330 -3961
rect -283 -3961 -249 -3943
rect -283 -3977 -249 -3961
rect -202 -3961 -168 -3943
rect -202 -3977 -168 -3961
rect -364 -4029 -330 -4015
rect -364 -4049 -330 -4029
rect -283 -4029 -249 -4015
rect -283 -4049 -249 -4029
rect -202 -4029 -168 -4015
rect -202 -4049 -168 -4029
rect -364 -4097 -330 -4087
rect -364 -4121 -330 -4097
rect -283 -4097 -249 -4087
rect -283 -4121 -249 -4097
rect -202 -4097 -168 -4087
rect -202 -4121 -168 -4097
rect -364 -4165 -330 -4159
rect -364 -4193 -330 -4165
rect -283 -4165 -249 -4159
rect -283 -4193 -249 -4165
rect -202 -4165 -168 -4159
rect -202 -4193 -168 -4165
rect -364 -4233 -330 -4231
rect -364 -4265 -330 -4233
rect -283 -4233 -249 -4231
rect -283 -4265 -249 -4233
rect -202 -4233 -168 -4231
rect -202 -4265 -168 -4233
rect -364 -4335 -330 -4303
rect -364 -4337 -330 -4335
rect -283 -4335 -249 -4303
rect -283 -4337 -249 -4335
rect -202 -4335 -168 -4303
rect -202 -4337 -168 -4335
rect -364 -4403 -330 -4375
rect -364 -4409 -330 -4403
rect -283 -4403 -249 -4375
rect -283 -4409 -249 -4403
rect -202 -4403 -168 -4375
rect -202 -4409 -168 -4403
rect -364 -4471 -330 -4447
rect -364 -4481 -330 -4471
rect -283 -4471 -249 -4447
rect -283 -4481 -249 -4471
rect -202 -4471 -168 -4447
rect -202 -4481 -168 -4471
rect -364 -4539 -330 -4519
rect -364 -4553 -330 -4539
rect -283 -4539 -249 -4519
rect -283 -4553 -249 -4539
rect -202 -4539 -168 -4519
rect -202 -4553 -168 -4539
rect -364 -4607 -330 -4591
rect -364 -4625 -330 -4607
rect -283 -4607 -249 -4591
rect -283 -4625 -249 -4607
rect -202 -4607 -168 -4591
rect -202 -4625 -168 -4607
rect -364 -4675 -330 -4663
rect -364 -4697 -330 -4675
rect -283 -4675 -249 -4663
rect -283 -4697 -249 -4675
rect -202 -4675 -168 -4663
rect -202 -4697 -168 -4675
rect -364 -4743 -330 -4735
rect -364 -4769 -330 -4743
rect -283 -4743 -249 -4735
rect -283 -4769 -249 -4743
rect -202 -4743 -168 -4735
rect -202 -4769 -168 -4743
rect -364 -4811 -330 -4807
rect -364 -4841 -330 -4811
rect -283 -4811 -249 -4807
rect -283 -4841 -249 -4811
rect -202 -4811 -168 -4807
rect -202 -4841 -168 -4811
rect -364 -4913 -330 -4879
rect -283 -4913 -249 -4879
rect -202 -4913 -168 -4879
rect -364 -4981 -330 -4951
rect -364 -4985 -330 -4981
rect -283 -4981 -249 -4951
rect -283 -4985 -249 -4981
rect -202 -4981 -168 -4951
rect -202 -4985 -168 -4981
rect -53 4981 53 4985
rect -53 -4981 53 4981
rect -53 -4985 53 -4981
rect 168 4981 202 4985
rect 168 4951 202 4981
rect 249 4981 283 4985
rect 249 4951 283 4981
rect 330 4981 364 4985
rect 330 4951 364 4981
rect 168 4879 202 4913
rect 249 4879 283 4913
rect 330 4879 364 4913
rect 168 4811 202 4841
rect 168 4807 202 4811
rect 249 4811 283 4841
rect 249 4807 283 4811
rect 330 4811 364 4841
rect 330 4807 364 4811
rect 168 4743 202 4769
rect 168 4735 202 4743
rect 249 4743 283 4769
rect 249 4735 283 4743
rect 330 4743 364 4769
rect 330 4735 364 4743
rect 168 4675 202 4697
rect 168 4663 202 4675
rect 249 4675 283 4697
rect 249 4663 283 4675
rect 330 4675 364 4697
rect 330 4663 364 4675
rect 168 4607 202 4625
rect 168 4591 202 4607
rect 249 4607 283 4625
rect 249 4591 283 4607
rect 330 4607 364 4625
rect 330 4591 364 4607
rect 168 4539 202 4553
rect 168 4519 202 4539
rect 249 4539 283 4553
rect 249 4519 283 4539
rect 330 4539 364 4553
rect 330 4519 364 4539
rect 168 4471 202 4481
rect 168 4447 202 4471
rect 249 4471 283 4481
rect 249 4447 283 4471
rect 330 4471 364 4481
rect 330 4447 364 4471
rect 168 4403 202 4409
rect 168 4375 202 4403
rect 249 4403 283 4409
rect 249 4375 283 4403
rect 330 4403 364 4409
rect 330 4375 364 4403
rect 168 4335 202 4337
rect 168 4303 202 4335
rect 249 4335 283 4337
rect 249 4303 283 4335
rect 330 4335 364 4337
rect 330 4303 364 4335
rect 168 4233 202 4265
rect 168 4231 202 4233
rect 249 4233 283 4265
rect 249 4231 283 4233
rect 330 4233 364 4265
rect 330 4231 364 4233
rect 168 4165 202 4193
rect 168 4159 202 4165
rect 249 4165 283 4193
rect 249 4159 283 4165
rect 330 4165 364 4193
rect 330 4159 364 4165
rect 168 4097 202 4121
rect 168 4087 202 4097
rect 249 4097 283 4121
rect 249 4087 283 4097
rect 330 4097 364 4121
rect 330 4087 364 4097
rect 168 4029 202 4049
rect 168 4015 202 4029
rect 249 4029 283 4049
rect 249 4015 283 4029
rect 330 4029 364 4049
rect 330 4015 364 4029
rect 168 3961 202 3977
rect 168 3943 202 3961
rect 249 3961 283 3977
rect 249 3943 283 3961
rect 330 3961 364 3977
rect 330 3943 364 3961
rect 168 3893 202 3905
rect 168 3871 202 3893
rect 249 3893 283 3905
rect 249 3871 283 3893
rect 330 3893 364 3905
rect 330 3871 364 3893
rect 168 3825 202 3833
rect 168 3799 202 3825
rect 249 3825 283 3833
rect 249 3799 283 3825
rect 330 3825 364 3833
rect 330 3799 364 3825
rect 168 3757 202 3761
rect 168 3727 202 3757
rect 249 3757 283 3761
rect 249 3727 283 3757
rect 330 3757 364 3761
rect 330 3727 364 3757
rect 168 3655 202 3689
rect 249 3655 283 3689
rect 330 3655 364 3689
rect 168 3587 202 3617
rect 168 3583 202 3587
rect 249 3587 283 3617
rect 249 3583 283 3587
rect 330 3587 364 3617
rect 330 3583 364 3587
rect 168 3519 202 3545
rect 168 3511 202 3519
rect 249 3519 283 3545
rect 249 3511 283 3519
rect 330 3519 364 3545
rect 330 3511 364 3519
rect 168 3451 202 3473
rect 168 3439 202 3451
rect 249 3451 283 3473
rect 249 3439 283 3451
rect 330 3451 364 3473
rect 330 3439 364 3451
rect 168 3383 202 3401
rect 168 3367 202 3383
rect 249 3383 283 3401
rect 249 3367 283 3383
rect 330 3383 364 3401
rect 330 3367 364 3383
rect 168 3315 202 3329
rect 168 3295 202 3315
rect 249 3315 283 3329
rect 249 3295 283 3315
rect 330 3315 364 3329
rect 330 3295 364 3315
rect 168 3247 202 3257
rect 168 3223 202 3247
rect 249 3247 283 3257
rect 249 3223 283 3247
rect 330 3247 364 3257
rect 330 3223 364 3247
rect 168 3179 202 3185
rect 168 3151 202 3179
rect 249 3179 283 3185
rect 249 3151 283 3179
rect 330 3179 364 3185
rect 330 3151 364 3179
rect 168 3111 202 3113
rect 168 3079 202 3111
rect 249 3111 283 3113
rect 249 3079 283 3111
rect 330 3111 364 3113
rect 330 3079 364 3111
rect 168 3009 202 3041
rect 168 3007 202 3009
rect 249 3009 283 3041
rect 249 3007 283 3009
rect 330 3009 364 3041
rect 330 3007 364 3009
rect 168 2941 202 2969
rect 168 2935 202 2941
rect 249 2941 283 2969
rect 249 2935 283 2941
rect 330 2941 364 2969
rect 330 2935 364 2941
rect 168 2873 202 2897
rect 168 2863 202 2873
rect 249 2873 283 2897
rect 249 2863 283 2873
rect 330 2873 364 2897
rect 330 2863 364 2873
rect 168 2805 202 2825
rect 168 2791 202 2805
rect 249 2805 283 2825
rect 249 2791 283 2805
rect 330 2805 364 2825
rect 330 2791 364 2805
rect 168 2737 202 2753
rect 168 2719 202 2737
rect 249 2737 283 2753
rect 249 2719 283 2737
rect 330 2737 364 2753
rect 330 2719 364 2737
rect 168 2669 202 2681
rect 168 2647 202 2669
rect 249 2669 283 2681
rect 249 2647 283 2669
rect 330 2669 364 2681
rect 330 2647 364 2669
rect 168 2601 202 2609
rect 168 2575 202 2601
rect 249 2601 283 2609
rect 249 2575 283 2601
rect 330 2601 364 2609
rect 330 2575 364 2601
rect 168 2533 202 2537
rect 168 2503 202 2533
rect 249 2533 283 2537
rect 249 2503 283 2533
rect 330 2533 364 2537
rect 330 2503 364 2533
rect 168 2431 202 2465
rect 249 2431 283 2465
rect 330 2431 364 2465
rect 168 2363 202 2393
rect 168 2359 202 2363
rect 249 2363 283 2393
rect 249 2359 283 2363
rect 330 2363 364 2393
rect 330 2359 364 2363
rect 168 2295 202 2321
rect 168 2287 202 2295
rect 249 2295 283 2321
rect 249 2287 283 2295
rect 330 2295 364 2321
rect 330 2287 364 2295
rect 168 2227 202 2249
rect 168 2215 202 2227
rect 249 2227 283 2249
rect 249 2215 283 2227
rect 330 2227 364 2249
rect 330 2215 364 2227
rect 168 2159 202 2177
rect 168 2143 202 2159
rect 249 2159 283 2177
rect 249 2143 283 2159
rect 330 2159 364 2177
rect 330 2143 364 2159
rect 168 2091 202 2105
rect 168 2071 202 2091
rect 249 2091 283 2105
rect 249 2071 283 2091
rect 330 2091 364 2105
rect 330 2071 364 2091
rect 168 2023 202 2033
rect 168 1999 202 2023
rect 249 2023 283 2033
rect 249 1999 283 2023
rect 330 2023 364 2033
rect 330 1999 364 2023
rect 168 1955 202 1961
rect 168 1927 202 1955
rect 249 1955 283 1961
rect 249 1927 283 1955
rect 330 1955 364 1961
rect 330 1927 364 1955
rect 168 1887 202 1889
rect 168 1855 202 1887
rect 249 1887 283 1889
rect 249 1855 283 1887
rect 330 1887 364 1889
rect 330 1855 364 1887
rect 168 1785 202 1817
rect 168 1783 202 1785
rect 249 1785 283 1817
rect 249 1783 283 1785
rect 330 1785 364 1817
rect 330 1783 364 1785
rect 168 1717 202 1745
rect 168 1711 202 1717
rect 249 1717 283 1745
rect 249 1711 283 1717
rect 330 1717 364 1745
rect 330 1711 364 1717
rect 168 1649 202 1673
rect 168 1639 202 1649
rect 249 1649 283 1673
rect 249 1639 283 1649
rect 330 1649 364 1673
rect 330 1639 364 1649
rect 168 1581 202 1601
rect 168 1567 202 1581
rect 249 1581 283 1601
rect 249 1567 283 1581
rect 330 1581 364 1601
rect 330 1567 364 1581
rect 168 1513 202 1529
rect 168 1495 202 1513
rect 249 1513 283 1529
rect 249 1495 283 1513
rect 330 1513 364 1529
rect 330 1495 364 1513
rect 168 1445 202 1457
rect 168 1423 202 1445
rect 249 1445 283 1457
rect 249 1423 283 1445
rect 330 1445 364 1457
rect 330 1423 364 1445
rect 168 1377 202 1385
rect 168 1351 202 1377
rect 249 1377 283 1385
rect 249 1351 283 1377
rect 330 1377 364 1385
rect 330 1351 364 1377
rect 168 1309 202 1313
rect 168 1279 202 1309
rect 249 1309 283 1313
rect 249 1279 283 1309
rect 330 1309 364 1313
rect 330 1279 364 1309
rect 168 1207 202 1241
rect 249 1207 283 1241
rect 330 1207 364 1241
rect 168 1139 202 1169
rect 168 1135 202 1139
rect 249 1139 283 1169
rect 249 1135 283 1139
rect 330 1139 364 1169
rect 330 1135 364 1139
rect 168 1071 202 1097
rect 168 1063 202 1071
rect 249 1071 283 1097
rect 249 1063 283 1071
rect 330 1071 364 1097
rect 330 1063 364 1071
rect 168 1003 202 1025
rect 168 991 202 1003
rect 249 1003 283 1025
rect 249 991 283 1003
rect 330 1003 364 1025
rect 330 991 364 1003
rect 168 935 202 953
rect 168 919 202 935
rect 249 935 283 953
rect 249 919 283 935
rect 330 935 364 953
rect 330 919 364 935
rect 168 867 202 881
rect 168 847 202 867
rect 249 867 283 881
rect 249 847 283 867
rect 330 867 364 881
rect 330 847 364 867
rect 168 799 202 809
rect 168 775 202 799
rect 249 799 283 809
rect 249 775 283 799
rect 330 799 364 809
rect 330 775 364 799
rect 168 731 202 737
rect 168 703 202 731
rect 249 731 283 737
rect 249 703 283 731
rect 330 731 364 737
rect 330 703 364 731
rect 168 663 202 665
rect 168 631 202 663
rect 249 663 283 665
rect 249 631 283 663
rect 330 663 364 665
rect 330 631 364 663
rect 168 561 202 593
rect 168 559 202 561
rect 249 561 283 593
rect 249 559 283 561
rect 330 561 364 593
rect 330 559 364 561
rect 168 493 202 521
rect 168 487 202 493
rect 249 493 283 521
rect 249 487 283 493
rect 330 493 364 521
rect 330 487 364 493
rect 168 425 202 449
rect 168 415 202 425
rect 249 425 283 449
rect 249 415 283 425
rect 330 425 364 449
rect 330 415 364 425
rect 168 357 202 377
rect 168 343 202 357
rect 249 357 283 377
rect 249 343 283 357
rect 330 357 364 377
rect 330 343 364 357
rect 168 289 202 305
rect 168 271 202 289
rect 249 289 283 305
rect 249 271 283 289
rect 330 289 364 305
rect 330 271 364 289
rect 168 221 202 233
rect 168 199 202 221
rect 249 221 283 233
rect 249 199 283 221
rect 330 221 364 233
rect 330 199 364 221
rect 168 153 202 161
rect 168 127 202 153
rect 249 153 283 161
rect 249 127 283 153
rect 330 153 364 161
rect 330 127 364 153
rect 168 85 202 89
rect 168 55 202 85
rect 249 85 283 89
rect 249 55 283 85
rect 330 85 364 89
rect 330 55 364 85
rect 168 -17 202 17
rect 249 -17 283 17
rect 330 -17 364 17
rect 168 -85 202 -55
rect 168 -89 202 -85
rect 249 -85 283 -55
rect 249 -89 283 -85
rect 330 -85 364 -55
rect 330 -89 364 -85
rect 168 -153 202 -127
rect 168 -161 202 -153
rect 249 -153 283 -127
rect 249 -161 283 -153
rect 330 -153 364 -127
rect 330 -161 364 -153
rect 168 -221 202 -199
rect 168 -233 202 -221
rect 249 -221 283 -199
rect 249 -233 283 -221
rect 330 -221 364 -199
rect 330 -233 364 -221
rect 168 -289 202 -271
rect 168 -305 202 -289
rect 249 -289 283 -271
rect 249 -305 283 -289
rect 330 -289 364 -271
rect 330 -305 364 -289
rect 168 -357 202 -343
rect 168 -377 202 -357
rect 249 -357 283 -343
rect 249 -377 283 -357
rect 330 -357 364 -343
rect 330 -377 364 -357
rect 168 -425 202 -415
rect 168 -449 202 -425
rect 249 -425 283 -415
rect 249 -449 283 -425
rect 330 -425 364 -415
rect 330 -449 364 -425
rect 168 -493 202 -487
rect 168 -521 202 -493
rect 249 -493 283 -487
rect 249 -521 283 -493
rect 330 -493 364 -487
rect 330 -521 364 -493
rect 168 -561 202 -559
rect 168 -593 202 -561
rect 249 -561 283 -559
rect 249 -593 283 -561
rect 330 -561 364 -559
rect 330 -593 364 -561
rect 168 -663 202 -631
rect 168 -665 202 -663
rect 249 -663 283 -631
rect 249 -665 283 -663
rect 330 -663 364 -631
rect 330 -665 364 -663
rect 168 -731 202 -703
rect 168 -737 202 -731
rect 249 -731 283 -703
rect 249 -737 283 -731
rect 330 -731 364 -703
rect 330 -737 364 -731
rect 168 -799 202 -775
rect 168 -809 202 -799
rect 249 -799 283 -775
rect 249 -809 283 -799
rect 330 -799 364 -775
rect 330 -809 364 -799
rect 168 -867 202 -847
rect 168 -881 202 -867
rect 249 -867 283 -847
rect 249 -881 283 -867
rect 330 -867 364 -847
rect 330 -881 364 -867
rect 168 -935 202 -919
rect 168 -953 202 -935
rect 249 -935 283 -919
rect 249 -953 283 -935
rect 330 -935 364 -919
rect 330 -953 364 -935
rect 168 -1003 202 -991
rect 168 -1025 202 -1003
rect 249 -1003 283 -991
rect 249 -1025 283 -1003
rect 330 -1003 364 -991
rect 330 -1025 364 -1003
rect 168 -1071 202 -1063
rect 168 -1097 202 -1071
rect 249 -1071 283 -1063
rect 249 -1097 283 -1071
rect 330 -1071 364 -1063
rect 330 -1097 364 -1071
rect 168 -1139 202 -1135
rect 168 -1169 202 -1139
rect 249 -1139 283 -1135
rect 249 -1169 283 -1139
rect 330 -1139 364 -1135
rect 330 -1169 364 -1139
rect 168 -1241 202 -1207
rect 249 -1241 283 -1207
rect 330 -1241 364 -1207
rect 168 -1309 202 -1279
rect 168 -1313 202 -1309
rect 249 -1309 283 -1279
rect 249 -1313 283 -1309
rect 330 -1309 364 -1279
rect 330 -1313 364 -1309
rect 168 -1377 202 -1351
rect 168 -1385 202 -1377
rect 249 -1377 283 -1351
rect 249 -1385 283 -1377
rect 330 -1377 364 -1351
rect 330 -1385 364 -1377
rect 168 -1445 202 -1423
rect 168 -1457 202 -1445
rect 249 -1445 283 -1423
rect 249 -1457 283 -1445
rect 330 -1445 364 -1423
rect 330 -1457 364 -1445
rect 168 -1513 202 -1495
rect 168 -1529 202 -1513
rect 249 -1513 283 -1495
rect 249 -1529 283 -1513
rect 330 -1513 364 -1495
rect 330 -1529 364 -1513
rect 168 -1581 202 -1567
rect 168 -1601 202 -1581
rect 249 -1581 283 -1567
rect 249 -1601 283 -1581
rect 330 -1581 364 -1567
rect 330 -1601 364 -1581
rect 168 -1649 202 -1639
rect 168 -1673 202 -1649
rect 249 -1649 283 -1639
rect 249 -1673 283 -1649
rect 330 -1649 364 -1639
rect 330 -1673 364 -1649
rect 168 -1717 202 -1711
rect 168 -1745 202 -1717
rect 249 -1717 283 -1711
rect 249 -1745 283 -1717
rect 330 -1717 364 -1711
rect 330 -1745 364 -1717
rect 168 -1785 202 -1783
rect 168 -1817 202 -1785
rect 249 -1785 283 -1783
rect 249 -1817 283 -1785
rect 330 -1785 364 -1783
rect 330 -1817 364 -1785
rect 168 -1887 202 -1855
rect 168 -1889 202 -1887
rect 249 -1887 283 -1855
rect 249 -1889 283 -1887
rect 330 -1887 364 -1855
rect 330 -1889 364 -1887
rect 168 -1955 202 -1927
rect 168 -1961 202 -1955
rect 249 -1955 283 -1927
rect 249 -1961 283 -1955
rect 330 -1955 364 -1927
rect 330 -1961 364 -1955
rect 168 -2023 202 -1999
rect 168 -2033 202 -2023
rect 249 -2023 283 -1999
rect 249 -2033 283 -2023
rect 330 -2023 364 -1999
rect 330 -2033 364 -2023
rect 168 -2091 202 -2071
rect 168 -2105 202 -2091
rect 249 -2091 283 -2071
rect 249 -2105 283 -2091
rect 330 -2091 364 -2071
rect 330 -2105 364 -2091
rect 168 -2159 202 -2143
rect 168 -2177 202 -2159
rect 249 -2159 283 -2143
rect 249 -2177 283 -2159
rect 330 -2159 364 -2143
rect 330 -2177 364 -2159
rect 168 -2227 202 -2215
rect 168 -2249 202 -2227
rect 249 -2227 283 -2215
rect 249 -2249 283 -2227
rect 330 -2227 364 -2215
rect 330 -2249 364 -2227
rect 168 -2295 202 -2287
rect 168 -2321 202 -2295
rect 249 -2295 283 -2287
rect 249 -2321 283 -2295
rect 330 -2295 364 -2287
rect 330 -2321 364 -2295
rect 168 -2363 202 -2359
rect 168 -2393 202 -2363
rect 249 -2363 283 -2359
rect 249 -2393 283 -2363
rect 330 -2363 364 -2359
rect 330 -2393 364 -2363
rect 168 -2465 202 -2431
rect 249 -2465 283 -2431
rect 330 -2465 364 -2431
rect 168 -2533 202 -2503
rect 168 -2537 202 -2533
rect 249 -2533 283 -2503
rect 249 -2537 283 -2533
rect 330 -2533 364 -2503
rect 330 -2537 364 -2533
rect 168 -2601 202 -2575
rect 168 -2609 202 -2601
rect 249 -2601 283 -2575
rect 249 -2609 283 -2601
rect 330 -2601 364 -2575
rect 330 -2609 364 -2601
rect 168 -2669 202 -2647
rect 168 -2681 202 -2669
rect 249 -2669 283 -2647
rect 249 -2681 283 -2669
rect 330 -2669 364 -2647
rect 330 -2681 364 -2669
rect 168 -2737 202 -2719
rect 168 -2753 202 -2737
rect 249 -2737 283 -2719
rect 249 -2753 283 -2737
rect 330 -2737 364 -2719
rect 330 -2753 364 -2737
rect 168 -2805 202 -2791
rect 168 -2825 202 -2805
rect 249 -2805 283 -2791
rect 249 -2825 283 -2805
rect 330 -2805 364 -2791
rect 330 -2825 364 -2805
rect 168 -2873 202 -2863
rect 168 -2897 202 -2873
rect 249 -2873 283 -2863
rect 249 -2897 283 -2873
rect 330 -2873 364 -2863
rect 330 -2897 364 -2873
rect 168 -2941 202 -2935
rect 168 -2969 202 -2941
rect 249 -2941 283 -2935
rect 249 -2969 283 -2941
rect 330 -2941 364 -2935
rect 330 -2969 364 -2941
rect 168 -3009 202 -3007
rect 168 -3041 202 -3009
rect 249 -3009 283 -3007
rect 249 -3041 283 -3009
rect 330 -3009 364 -3007
rect 330 -3041 364 -3009
rect 168 -3111 202 -3079
rect 168 -3113 202 -3111
rect 249 -3111 283 -3079
rect 249 -3113 283 -3111
rect 330 -3111 364 -3079
rect 330 -3113 364 -3111
rect 168 -3179 202 -3151
rect 168 -3185 202 -3179
rect 249 -3179 283 -3151
rect 249 -3185 283 -3179
rect 330 -3179 364 -3151
rect 330 -3185 364 -3179
rect 168 -3247 202 -3223
rect 168 -3257 202 -3247
rect 249 -3247 283 -3223
rect 249 -3257 283 -3247
rect 330 -3247 364 -3223
rect 330 -3257 364 -3247
rect 168 -3315 202 -3295
rect 168 -3329 202 -3315
rect 249 -3315 283 -3295
rect 249 -3329 283 -3315
rect 330 -3315 364 -3295
rect 330 -3329 364 -3315
rect 168 -3383 202 -3367
rect 168 -3401 202 -3383
rect 249 -3383 283 -3367
rect 249 -3401 283 -3383
rect 330 -3383 364 -3367
rect 330 -3401 364 -3383
rect 168 -3451 202 -3439
rect 168 -3473 202 -3451
rect 249 -3451 283 -3439
rect 249 -3473 283 -3451
rect 330 -3451 364 -3439
rect 330 -3473 364 -3451
rect 168 -3519 202 -3511
rect 168 -3545 202 -3519
rect 249 -3519 283 -3511
rect 249 -3545 283 -3519
rect 330 -3519 364 -3511
rect 330 -3545 364 -3519
rect 168 -3587 202 -3583
rect 168 -3617 202 -3587
rect 249 -3587 283 -3583
rect 249 -3617 283 -3587
rect 330 -3587 364 -3583
rect 330 -3617 364 -3587
rect 168 -3689 202 -3655
rect 249 -3689 283 -3655
rect 330 -3689 364 -3655
rect 168 -3757 202 -3727
rect 168 -3761 202 -3757
rect 249 -3757 283 -3727
rect 249 -3761 283 -3757
rect 330 -3757 364 -3727
rect 330 -3761 364 -3757
rect 168 -3825 202 -3799
rect 168 -3833 202 -3825
rect 249 -3825 283 -3799
rect 249 -3833 283 -3825
rect 330 -3825 364 -3799
rect 330 -3833 364 -3825
rect 168 -3893 202 -3871
rect 168 -3905 202 -3893
rect 249 -3893 283 -3871
rect 249 -3905 283 -3893
rect 330 -3893 364 -3871
rect 330 -3905 364 -3893
rect 168 -3961 202 -3943
rect 168 -3977 202 -3961
rect 249 -3961 283 -3943
rect 249 -3977 283 -3961
rect 330 -3961 364 -3943
rect 330 -3977 364 -3961
rect 168 -4029 202 -4015
rect 168 -4049 202 -4029
rect 249 -4029 283 -4015
rect 249 -4049 283 -4029
rect 330 -4029 364 -4015
rect 330 -4049 364 -4029
rect 168 -4097 202 -4087
rect 168 -4121 202 -4097
rect 249 -4097 283 -4087
rect 249 -4121 283 -4097
rect 330 -4097 364 -4087
rect 330 -4121 364 -4097
rect 168 -4165 202 -4159
rect 168 -4193 202 -4165
rect 249 -4165 283 -4159
rect 249 -4193 283 -4165
rect 330 -4165 364 -4159
rect 330 -4193 364 -4165
rect 168 -4233 202 -4231
rect 168 -4265 202 -4233
rect 249 -4233 283 -4231
rect 249 -4265 283 -4233
rect 330 -4233 364 -4231
rect 330 -4265 364 -4233
rect 168 -4335 202 -4303
rect 168 -4337 202 -4335
rect 249 -4335 283 -4303
rect 249 -4337 283 -4335
rect 330 -4335 364 -4303
rect 330 -4337 364 -4335
rect 168 -4403 202 -4375
rect 168 -4409 202 -4403
rect 249 -4403 283 -4375
rect 249 -4409 283 -4403
rect 330 -4403 364 -4375
rect 330 -4409 364 -4403
rect 168 -4471 202 -4447
rect 168 -4481 202 -4471
rect 249 -4471 283 -4447
rect 249 -4481 283 -4471
rect 330 -4471 364 -4447
rect 330 -4481 364 -4471
rect 168 -4539 202 -4519
rect 168 -4553 202 -4539
rect 249 -4539 283 -4519
rect 249 -4553 283 -4539
rect 330 -4539 364 -4519
rect 330 -4553 364 -4539
rect 168 -4607 202 -4591
rect 168 -4625 202 -4607
rect 249 -4607 283 -4591
rect 249 -4625 283 -4607
rect 330 -4607 364 -4591
rect 330 -4625 364 -4607
rect 168 -4675 202 -4663
rect 168 -4697 202 -4675
rect 249 -4675 283 -4663
rect 249 -4697 283 -4675
rect 330 -4675 364 -4663
rect 330 -4697 364 -4675
rect 168 -4743 202 -4735
rect 168 -4769 202 -4743
rect 249 -4743 283 -4735
rect 249 -4769 283 -4743
rect 330 -4743 364 -4735
rect 330 -4769 364 -4743
rect 168 -4811 202 -4807
rect 168 -4841 202 -4811
rect 249 -4811 283 -4807
rect 249 -4841 283 -4811
rect 330 -4811 364 -4807
rect 330 -4841 364 -4811
rect 168 -4913 202 -4879
rect 249 -4913 283 -4879
rect 330 -4913 364 -4879
rect 168 -4981 202 -4951
rect 168 -4985 202 -4981
rect 249 -4981 283 -4951
rect 249 -4985 283 -4981
rect 330 -4981 364 -4951
rect 330 -4985 364 -4981
rect 479 4981 585 4985
rect 479 -4981 585 4981
rect 479 -4985 585 -4981
rect 700 4981 734 4985
rect 700 4951 734 4981
rect 781 4981 815 4985
rect 781 4951 815 4981
rect 862 4981 896 4985
rect 862 4951 896 4981
rect 700 4879 734 4913
rect 781 4879 815 4913
rect 862 4879 896 4913
rect 700 4811 734 4841
rect 700 4807 734 4811
rect 781 4811 815 4841
rect 781 4807 815 4811
rect 862 4811 896 4841
rect 862 4807 896 4811
rect 700 4743 734 4769
rect 700 4735 734 4743
rect 781 4743 815 4769
rect 781 4735 815 4743
rect 862 4743 896 4769
rect 862 4735 896 4743
rect 700 4675 734 4697
rect 700 4663 734 4675
rect 781 4675 815 4697
rect 781 4663 815 4675
rect 862 4675 896 4697
rect 862 4663 896 4675
rect 700 4607 734 4625
rect 700 4591 734 4607
rect 781 4607 815 4625
rect 781 4591 815 4607
rect 862 4607 896 4625
rect 862 4591 896 4607
rect 700 4539 734 4553
rect 700 4519 734 4539
rect 781 4539 815 4553
rect 781 4519 815 4539
rect 862 4539 896 4553
rect 862 4519 896 4539
rect 700 4471 734 4481
rect 700 4447 734 4471
rect 781 4471 815 4481
rect 781 4447 815 4471
rect 862 4471 896 4481
rect 862 4447 896 4471
rect 700 4403 734 4409
rect 700 4375 734 4403
rect 781 4403 815 4409
rect 781 4375 815 4403
rect 862 4403 896 4409
rect 862 4375 896 4403
rect 700 4335 734 4337
rect 700 4303 734 4335
rect 781 4335 815 4337
rect 781 4303 815 4335
rect 862 4335 896 4337
rect 862 4303 896 4335
rect 700 4233 734 4265
rect 700 4231 734 4233
rect 781 4233 815 4265
rect 781 4231 815 4233
rect 862 4233 896 4265
rect 862 4231 896 4233
rect 700 4165 734 4193
rect 700 4159 734 4165
rect 781 4165 815 4193
rect 781 4159 815 4165
rect 862 4165 896 4193
rect 862 4159 896 4165
rect 700 4097 734 4121
rect 700 4087 734 4097
rect 781 4097 815 4121
rect 781 4087 815 4097
rect 862 4097 896 4121
rect 862 4087 896 4097
rect 700 4029 734 4049
rect 700 4015 734 4029
rect 781 4029 815 4049
rect 781 4015 815 4029
rect 862 4029 896 4049
rect 862 4015 896 4029
rect 700 3961 734 3977
rect 700 3943 734 3961
rect 781 3961 815 3977
rect 781 3943 815 3961
rect 862 3961 896 3977
rect 862 3943 896 3961
rect 700 3893 734 3905
rect 700 3871 734 3893
rect 781 3893 815 3905
rect 781 3871 815 3893
rect 862 3893 896 3905
rect 862 3871 896 3893
rect 700 3825 734 3833
rect 700 3799 734 3825
rect 781 3825 815 3833
rect 781 3799 815 3825
rect 862 3825 896 3833
rect 862 3799 896 3825
rect 700 3757 734 3761
rect 700 3727 734 3757
rect 781 3757 815 3761
rect 781 3727 815 3757
rect 862 3757 896 3761
rect 862 3727 896 3757
rect 700 3655 734 3689
rect 781 3655 815 3689
rect 862 3655 896 3689
rect 700 3587 734 3617
rect 700 3583 734 3587
rect 781 3587 815 3617
rect 781 3583 815 3587
rect 862 3587 896 3617
rect 862 3583 896 3587
rect 700 3519 734 3545
rect 700 3511 734 3519
rect 781 3519 815 3545
rect 781 3511 815 3519
rect 862 3519 896 3545
rect 862 3511 896 3519
rect 700 3451 734 3473
rect 700 3439 734 3451
rect 781 3451 815 3473
rect 781 3439 815 3451
rect 862 3451 896 3473
rect 862 3439 896 3451
rect 700 3383 734 3401
rect 700 3367 734 3383
rect 781 3383 815 3401
rect 781 3367 815 3383
rect 862 3383 896 3401
rect 862 3367 896 3383
rect 700 3315 734 3329
rect 700 3295 734 3315
rect 781 3315 815 3329
rect 781 3295 815 3315
rect 862 3315 896 3329
rect 862 3295 896 3315
rect 700 3247 734 3257
rect 700 3223 734 3247
rect 781 3247 815 3257
rect 781 3223 815 3247
rect 862 3247 896 3257
rect 862 3223 896 3247
rect 700 3179 734 3185
rect 700 3151 734 3179
rect 781 3179 815 3185
rect 781 3151 815 3179
rect 862 3179 896 3185
rect 862 3151 896 3179
rect 700 3111 734 3113
rect 700 3079 734 3111
rect 781 3111 815 3113
rect 781 3079 815 3111
rect 862 3111 896 3113
rect 862 3079 896 3111
rect 700 3009 734 3041
rect 700 3007 734 3009
rect 781 3009 815 3041
rect 781 3007 815 3009
rect 862 3009 896 3041
rect 862 3007 896 3009
rect 700 2941 734 2969
rect 700 2935 734 2941
rect 781 2941 815 2969
rect 781 2935 815 2941
rect 862 2941 896 2969
rect 862 2935 896 2941
rect 700 2873 734 2897
rect 700 2863 734 2873
rect 781 2873 815 2897
rect 781 2863 815 2873
rect 862 2873 896 2897
rect 862 2863 896 2873
rect 700 2805 734 2825
rect 700 2791 734 2805
rect 781 2805 815 2825
rect 781 2791 815 2805
rect 862 2805 896 2825
rect 862 2791 896 2805
rect 700 2737 734 2753
rect 700 2719 734 2737
rect 781 2737 815 2753
rect 781 2719 815 2737
rect 862 2737 896 2753
rect 862 2719 896 2737
rect 700 2669 734 2681
rect 700 2647 734 2669
rect 781 2669 815 2681
rect 781 2647 815 2669
rect 862 2669 896 2681
rect 862 2647 896 2669
rect 700 2601 734 2609
rect 700 2575 734 2601
rect 781 2601 815 2609
rect 781 2575 815 2601
rect 862 2601 896 2609
rect 862 2575 896 2601
rect 700 2533 734 2537
rect 700 2503 734 2533
rect 781 2533 815 2537
rect 781 2503 815 2533
rect 862 2533 896 2537
rect 862 2503 896 2533
rect 700 2431 734 2465
rect 781 2431 815 2465
rect 862 2431 896 2465
rect 700 2363 734 2393
rect 700 2359 734 2363
rect 781 2363 815 2393
rect 781 2359 815 2363
rect 862 2363 896 2393
rect 862 2359 896 2363
rect 700 2295 734 2321
rect 700 2287 734 2295
rect 781 2295 815 2321
rect 781 2287 815 2295
rect 862 2295 896 2321
rect 862 2287 896 2295
rect 700 2227 734 2249
rect 700 2215 734 2227
rect 781 2227 815 2249
rect 781 2215 815 2227
rect 862 2227 896 2249
rect 862 2215 896 2227
rect 700 2159 734 2177
rect 700 2143 734 2159
rect 781 2159 815 2177
rect 781 2143 815 2159
rect 862 2159 896 2177
rect 862 2143 896 2159
rect 700 2091 734 2105
rect 700 2071 734 2091
rect 781 2091 815 2105
rect 781 2071 815 2091
rect 862 2091 896 2105
rect 862 2071 896 2091
rect 700 2023 734 2033
rect 700 1999 734 2023
rect 781 2023 815 2033
rect 781 1999 815 2023
rect 862 2023 896 2033
rect 862 1999 896 2023
rect 700 1955 734 1961
rect 700 1927 734 1955
rect 781 1955 815 1961
rect 781 1927 815 1955
rect 862 1955 896 1961
rect 862 1927 896 1955
rect 700 1887 734 1889
rect 700 1855 734 1887
rect 781 1887 815 1889
rect 781 1855 815 1887
rect 862 1887 896 1889
rect 862 1855 896 1887
rect 700 1785 734 1817
rect 700 1783 734 1785
rect 781 1785 815 1817
rect 781 1783 815 1785
rect 862 1785 896 1817
rect 862 1783 896 1785
rect 700 1717 734 1745
rect 700 1711 734 1717
rect 781 1717 815 1745
rect 781 1711 815 1717
rect 862 1717 896 1745
rect 862 1711 896 1717
rect 700 1649 734 1673
rect 700 1639 734 1649
rect 781 1649 815 1673
rect 781 1639 815 1649
rect 862 1649 896 1673
rect 862 1639 896 1649
rect 700 1581 734 1601
rect 700 1567 734 1581
rect 781 1581 815 1601
rect 781 1567 815 1581
rect 862 1581 896 1601
rect 862 1567 896 1581
rect 700 1513 734 1529
rect 700 1495 734 1513
rect 781 1513 815 1529
rect 781 1495 815 1513
rect 862 1513 896 1529
rect 862 1495 896 1513
rect 700 1445 734 1457
rect 700 1423 734 1445
rect 781 1445 815 1457
rect 781 1423 815 1445
rect 862 1445 896 1457
rect 862 1423 896 1445
rect 700 1377 734 1385
rect 700 1351 734 1377
rect 781 1377 815 1385
rect 781 1351 815 1377
rect 862 1377 896 1385
rect 862 1351 896 1377
rect 700 1309 734 1313
rect 700 1279 734 1309
rect 781 1309 815 1313
rect 781 1279 815 1309
rect 862 1309 896 1313
rect 862 1279 896 1309
rect 700 1207 734 1241
rect 781 1207 815 1241
rect 862 1207 896 1241
rect 700 1139 734 1169
rect 700 1135 734 1139
rect 781 1139 815 1169
rect 781 1135 815 1139
rect 862 1139 896 1169
rect 862 1135 896 1139
rect 700 1071 734 1097
rect 700 1063 734 1071
rect 781 1071 815 1097
rect 781 1063 815 1071
rect 862 1071 896 1097
rect 862 1063 896 1071
rect 700 1003 734 1025
rect 700 991 734 1003
rect 781 1003 815 1025
rect 781 991 815 1003
rect 862 1003 896 1025
rect 862 991 896 1003
rect 700 935 734 953
rect 700 919 734 935
rect 781 935 815 953
rect 781 919 815 935
rect 862 935 896 953
rect 862 919 896 935
rect 700 867 734 881
rect 700 847 734 867
rect 781 867 815 881
rect 781 847 815 867
rect 862 867 896 881
rect 862 847 896 867
rect 700 799 734 809
rect 700 775 734 799
rect 781 799 815 809
rect 781 775 815 799
rect 862 799 896 809
rect 862 775 896 799
rect 700 731 734 737
rect 700 703 734 731
rect 781 731 815 737
rect 781 703 815 731
rect 862 731 896 737
rect 862 703 896 731
rect 700 663 734 665
rect 700 631 734 663
rect 781 663 815 665
rect 781 631 815 663
rect 862 663 896 665
rect 862 631 896 663
rect 700 561 734 593
rect 700 559 734 561
rect 781 561 815 593
rect 781 559 815 561
rect 862 561 896 593
rect 862 559 896 561
rect 700 493 734 521
rect 700 487 734 493
rect 781 493 815 521
rect 781 487 815 493
rect 862 493 896 521
rect 862 487 896 493
rect 700 425 734 449
rect 700 415 734 425
rect 781 425 815 449
rect 781 415 815 425
rect 862 425 896 449
rect 862 415 896 425
rect 700 357 734 377
rect 700 343 734 357
rect 781 357 815 377
rect 781 343 815 357
rect 862 357 896 377
rect 862 343 896 357
rect 700 289 734 305
rect 700 271 734 289
rect 781 289 815 305
rect 781 271 815 289
rect 862 289 896 305
rect 862 271 896 289
rect 700 221 734 233
rect 700 199 734 221
rect 781 221 815 233
rect 781 199 815 221
rect 862 221 896 233
rect 862 199 896 221
rect 700 153 734 161
rect 700 127 734 153
rect 781 153 815 161
rect 781 127 815 153
rect 862 153 896 161
rect 862 127 896 153
rect 700 85 734 89
rect 700 55 734 85
rect 781 85 815 89
rect 781 55 815 85
rect 862 85 896 89
rect 862 55 896 85
rect 700 -17 734 17
rect 781 -17 815 17
rect 862 -17 896 17
rect 700 -85 734 -55
rect 700 -89 734 -85
rect 781 -85 815 -55
rect 781 -89 815 -85
rect 862 -85 896 -55
rect 862 -89 896 -85
rect 700 -153 734 -127
rect 700 -161 734 -153
rect 781 -153 815 -127
rect 781 -161 815 -153
rect 862 -153 896 -127
rect 862 -161 896 -153
rect 700 -221 734 -199
rect 700 -233 734 -221
rect 781 -221 815 -199
rect 781 -233 815 -221
rect 862 -221 896 -199
rect 862 -233 896 -221
rect 700 -289 734 -271
rect 700 -305 734 -289
rect 781 -289 815 -271
rect 781 -305 815 -289
rect 862 -289 896 -271
rect 862 -305 896 -289
rect 700 -357 734 -343
rect 700 -377 734 -357
rect 781 -357 815 -343
rect 781 -377 815 -357
rect 862 -357 896 -343
rect 862 -377 896 -357
rect 700 -425 734 -415
rect 700 -449 734 -425
rect 781 -425 815 -415
rect 781 -449 815 -425
rect 862 -425 896 -415
rect 862 -449 896 -425
rect 700 -493 734 -487
rect 700 -521 734 -493
rect 781 -493 815 -487
rect 781 -521 815 -493
rect 862 -493 896 -487
rect 862 -521 896 -493
rect 700 -561 734 -559
rect 700 -593 734 -561
rect 781 -561 815 -559
rect 781 -593 815 -561
rect 862 -561 896 -559
rect 862 -593 896 -561
rect 700 -663 734 -631
rect 700 -665 734 -663
rect 781 -663 815 -631
rect 781 -665 815 -663
rect 862 -663 896 -631
rect 862 -665 896 -663
rect 700 -731 734 -703
rect 700 -737 734 -731
rect 781 -731 815 -703
rect 781 -737 815 -731
rect 862 -731 896 -703
rect 862 -737 896 -731
rect 700 -799 734 -775
rect 700 -809 734 -799
rect 781 -799 815 -775
rect 781 -809 815 -799
rect 862 -799 896 -775
rect 862 -809 896 -799
rect 700 -867 734 -847
rect 700 -881 734 -867
rect 781 -867 815 -847
rect 781 -881 815 -867
rect 862 -867 896 -847
rect 862 -881 896 -867
rect 700 -935 734 -919
rect 700 -953 734 -935
rect 781 -935 815 -919
rect 781 -953 815 -935
rect 862 -935 896 -919
rect 862 -953 896 -935
rect 700 -1003 734 -991
rect 700 -1025 734 -1003
rect 781 -1003 815 -991
rect 781 -1025 815 -1003
rect 862 -1003 896 -991
rect 862 -1025 896 -1003
rect 700 -1071 734 -1063
rect 700 -1097 734 -1071
rect 781 -1071 815 -1063
rect 781 -1097 815 -1071
rect 862 -1071 896 -1063
rect 862 -1097 896 -1071
rect 700 -1139 734 -1135
rect 700 -1169 734 -1139
rect 781 -1139 815 -1135
rect 781 -1169 815 -1139
rect 862 -1139 896 -1135
rect 862 -1169 896 -1139
rect 700 -1241 734 -1207
rect 781 -1241 815 -1207
rect 862 -1241 896 -1207
rect 700 -1309 734 -1279
rect 700 -1313 734 -1309
rect 781 -1309 815 -1279
rect 781 -1313 815 -1309
rect 862 -1309 896 -1279
rect 862 -1313 896 -1309
rect 700 -1377 734 -1351
rect 700 -1385 734 -1377
rect 781 -1377 815 -1351
rect 781 -1385 815 -1377
rect 862 -1377 896 -1351
rect 862 -1385 896 -1377
rect 700 -1445 734 -1423
rect 700 -1457 734 -1445
rect 781 -1445 815 -1423
rect 781 -1457 815 -1445
rect 862 -1445 896 -1423
rect 862 -1457 896 -1445
rect 700 -1513 734 -1495
rect 700 -1529 734 -1513
rect 781 -1513 815 -1495
rect 781 -1529 815 -1513
rect 862 -1513 896 -1495
rect 862 -1529 896 -1513
rect 700 -1581 734 -1567
rect 700 -1601 734 -1581
rect 781 -1581 815 -1567
rect 781 -1601 815 -1581
rect 862 -1581 896 -1567
rect 862 -1601 896 -1581
rect 700 -1649 734 -1639
rect 700 -1673 734 -1649
rect 781 -1649 815 -1639
rect 781 -1673 815 -1649
rect 862 -1649 896 -1639
rect 862 -1673 896 -1649
rect 700 -1717 734 -1711
rect 700 -1745 734 -1717
rect 781 -1717 815 -1711
rect 781 -1745 815 -1717
rect 862 -1717 896 -1711
rect 862 -1745 896 -1717
rect 700 -1785 734 -1783
rect 700 -1817 734 -1785
rect 781 -1785 815 -1783
rect 781 -1817 815 -1785
rect 862 -1785 896 -1783
rect 862 -1817 896 -1785
rect 700 -1887 734 -1855
rect 700 -1889 734 -1887
rect 781 -1887 815 -1855
rect 781 -1889 815 -1887
rect 862 -1887 896 -1855
rect 862 -1889 896 -1887
rect 700 -1955 734 -1927
rect 700 -1961 734 -1955
rect 781 -1955 815 -1927
rect 781 -1961 815 -1955
rect 862 -1955 896 -1927
rect 862 -1961 896 -1955
rect 700 -2023 734 -1999
rect 700 -2033 734 -2023
rect 781 -2023 815 -1999
rect 781 -2033 815 -2023
rect 862 -2023 896 -1999
rect 862 -2033 896 -2023
rect 700 -2091 734 -2071
rect 700 -2105 734 -2091
rect 781 -2091 815 -2071
rect 781 -2105 815 -2091
rect 862 -2091 896 -2071
rect 862 -2105 896 -2091
rect 700 -2159 734 -2143
rect 700 -2177 734 -2159
rect 781 -2159 815 -2143
rect 781 -2177 815 -2159
rect 862 -2159 896 -2143
rect 862 -2177 896 -2159
rect 700 -2227 734 -2215
rect 700 -2249 734 -2227
rect 781 -2227 815 -2215
rect 781 -2249 815 -2227
rect 862 -2227 896 -2215
rect 862 -2249 896 -2227
rect 700 -2295 734 -2287
rect 700 -2321 734 -2295
rect 781 -2295 815 -2287
rect 781 -2321 815 -2295
rect 862 -2295 896 -2287
rect 862 -2321 896 -2295
rect 700 -2363 734 -2359
rect 700 -2393 734 -2363
rect 781 -2363 815 -2359
rect 781 -2393 815 -2363
rect 862 -2363 896 -2359
rect 862 -2393 896 -2363
rect 700 -2465 734 -2431
rect 781 -2465 815 -2431
rect 862 -2465 896 -2431
rect 700 -2533 734 -2503
rect 700 -2537 734 -2533
rect 781 -2533 815 -2503
rect 781 -2537 815 -2533
rect 862 -2533 896 -2503
rect 862 -2537 896 -2533
rect 700 -2601 734 -2575
rect 700 -2609 734 -2601
rect 781 -2601 815 -2575
rect 781 -2609 815 -2601
rect 862 -2601 896 -2575
rect 862 -2609 896 -2601
rect 700 -2669 734 -2647
rect 700 -2681 734 -2669
rect 781 -2669 815 -2647
rect 781 -2681 815 -2669
rect 862 -2669 896 -2647
rect 862 -2681 896 -2669
rect 700 -2737 734 -2719
rect 700 -2753 734 -2737
rect 781 -2737 815 -2719
rect 781 -2753 815 -2737
rect 862 -2737 896 -2719
rect 862 -2753 896 -2737
rect 700 -2805 734 -2791
rect 700 -2825 734 -2805
rect 781 -2805 815 -2791
rect 781 -2825 815 -2805
rect 862 -2805 896 -2791
rect 862 -2825 896 -2805
rect 700 -2873 734 -2863
rect 700 -2897 734 -2873
rect 781 -2873 815 -2863
rect 781 -2897 815 -2873
rect 862 -2873 896 -2863
rect 862 -2897 896 -2873
rect 700 -2941 734 -2935
rect 700 -2969 734 -2941
rect 781 -2941 815 -2935
rect 781 -2969 815 -2941
rect 862 -2941 896 -2935
rect 862 -2969 896 -2941
rect 700 -3009 734 -3007
rect 700 -3041 734 -3009
rect 781 -3009 815 -3007
rect 781 -3041 815 -3009
rect 862 -3009 896 -3007
rect 862 -3041 896 -3009
rect 700 -3111 734 -3079
rect 700 -3113 734 -3111
rect 781 -3111 815 -3079
rect 781 -3113 815 -3111
rect 862 -3111 896 -3079
rect 862 -3113 896 -3111
rect 700 -3179 734 -3151
rect 700 -3185 734 -3179
rect 781 -3179 815 -3151
rect 781 -3185 815 -3179
rect 862 -3179 896 -3151
rect 862 -3185 896 -3179
rect 700 -3247 734 -3223
rect 700 -3257 734 -3247
rect 781 -3247 815 -3223
rect 781 -3257 815 -3247
rect 862 -3247 896 -3223
rect 862 -3257 896 -3247
rect 700 -3315 734 -3295
rect 700 -3329 734 -3315
rect 781 -3315 815 -3295
rect 781 -3329 815 -3315
rect 862 -3315 896 -3295
rect 862 -3329 896 -3315
rect 700 -3383 734 -3367
rect 700 -3401 734 -3383
rect 781 -3383 815 -3367
rect 781 -3401 815 -3383
rect 862 -3383 896 -3367
rect 862 -3401 896 -3383
rect 700 -3451 734 -3439
rect 700 -3473 734 -3451
rect 781 -3451 815 -3439
rect 781 -3473 815 -3451
rect 862 -3451 896 -3439
rect 862 -3473 896 -3451
rect 700 -3519 734 -3511
rect 700 -3545 734 -3519
rect 781 -3519 815 -3511
rect 781 -3545 815 -3519
rect 862 -3519 896 -3511
rect 862 -3545 896 -3519
rect 700 -3587 734 -3583
rect 700 -3617 734 -3587
rect 781 -3587 815 -3583
rect 781 -3617 815 -3587
rect 862 -3587 896 -3583
rect 862 -3617 896 -3587
rect 700 -3689 734 -3655
rect 781 -3689 815 -3655
rect 862 -3689 896 -3655
rect 700 -3757 734 -3727
rect 700 -3761 734 -3757
rect 781 -3757 815 -3727
rect 781 -3761 815 -3757
rect 862 -3757 896 -3727
rect 862 -3761 896 -3757
rect 700 -3825 734 -3799
rect 700 -3833 734 -3825
rect 781 -3825 815 -3799
rect 781 -3833 815 -3825
rect 862 -3825 896 -3799
rect 862 -3833 896 -3825
rect 700 -3893 734 -3871
rect 700 -3905 734 -3893
rect 781 -3893 815 -3871
rect 781 -3905 815 -3893
rect 862 -3893 896 -3871
rect 862 -3905 896 -3893
rect 700 -3961 734 -3943
rect 700 -3977 734 -3961
rect 781 -3961 815 -3943
rect 781 -3977 815 -3961
rect 862 -3961 896 -3943
rect 862 -3977 896 -3961
rect 700 -4029 734 -4015
rect 700 -4049 734 -4029
rect 781 -4029 815 -4015
rect 781 -4049 815 -4029
rect 862 -4029 896 -4015
rect 862 -4049 896 -4029
rect 700 -4097 734 -4087
rect 700 -4121 734 -4097
rect 781 -4097 815 -4087
rect 781 -4121 815 -4097
rect 862 -4097 896 -4087
rect 862 -4121 896 -4097
rect 700 -4165 734 -4159
rect 700 -4193 734 -4165
rect 781 -4165 815 -4159
rect 781 -4193 815 -4165
rect 862 -4165 896 -4159
rect 862 -4193 896 -4165
rect 700 -4233 734 -4231
rect 700 -4265 734 -4233
rect 781 -4233 815 -4231
rect 781 -4265 815 -4233
rect 862 -4233 896 -4231
rect 862 -4265 896 -4233
rect 700 -4335 734 -4303
rect 700 -4337 734 -4335
rect 781 -4335 815 -4303
rect 781 -4337 815 -4335
rect 862 -4335 896 -4303
rect 862 -4337 896 -4335
rect 700 -4403 734 -4375
rect 700 -4409 734 -4403
rect 781 -4403 815 -4375
rect 781 -4409 815 -4403
rect 862 -4403 896 -4375
rect 862 -4409 896 -4403
rect 700 -4471 734 -4447
rect 700 -4481 734 -4471
rect 781 -4471 815 -4447
rect 781 -4481 815 -4471
rect 862 -4471 896 -4447
rect 862 -4481 896 -4471
rect 700 -4539 734 -4519
rect 700 -4553 734 -4539
rect 781 -4539 815 -4519
rect 781 -4553 815 -4539
rect 862 -4539 896 -4519
rect 862 -4553 896 -4539
rect 700 -4607 734 -4591
rect 700 -4625 734 -4607
rect 781 -4607 815 -4591
rect 781 -4625 815 -4607
rect 862 -4607 896 -4591
rect 862 -4625 896 -4607
rect 700 -4675 734 -4663
rect 700 -4697 734 -4675
rect 781 -4675 815 -4663
rect 781 -4697 815 -4675
rect 862 -4675 896 -4663
rect 862 -4697 896 -4675
rect 700 -4743 734 -4735
rect 700 -4769 734 -4743
rect 781 -4743 815 -4735
rect 781 -4769 815 -4743
rect 862 -4743 896 -4735
rect 862 -4769 896 -4743
rect 700 -4811 734 -4807
rect 700 -4841 734 -4811
rect 781 -4811 815 -4807
rect 781 -4841 815 -4811
rect 862 -4811 896 -4807
rect 862 -4841 896 -4811
rect 700 -4913 734 -4879
rect 781 -4913 815 -4879
rect 862 -4913 896 -4879
rect 700 -4981 734 -4951
rect 700 -4985 734 -4981
rect 781 -4981 815 -4951
rect 781 -4985 815 -4981
rect 862 -4981 896 -4951
rect 862 -4985 896 -4981
rect 1011 4981 1117 4985
rect 1011 -4981 1117 4981
rect 1011 -4985 1117 -4981
rect 1232 4981 1266 4985
rect 1232 4951 1266 4981
rect 1232 4879 1266 4913
rect 1232 4811 1266 4841
rect 1232 4807 1266 4811
rect 1232 4743 1266 4769
rect 1232 4735 1266 4743
rect 1232 4675 1266 4697
rect 1232 4663 1266 4675
rect 1232 4607 1266 4625
rect 1232 4591 1266 4607
rect 1232 4539 1266 4553
rect 1232 4519 1266 4539
rect 1232 4471 1266 4481
rect 1232 4447 1266 4471
rect 1232 4403 1266 4409
rect 1232 4375 1266 4403
rect 1232 4335 1266 4337
rect 1232 4303 1266 4335
rect 1232 4233 1266 4265
rect 1232 4231 1266 4233
rect 1232 4165 1266 4193
rect 1232 4159 1266 4165
rect 1232 4097 1266 4121
rect 1232 4087 1266 4097
rect 1232 4029 1266 4049
rect 1232 4015 1266 4029
rect 1232 3961 1266 3977
rect 1232 3943 1266 3961
rect 1232 3893 1266 3905
rect 1232 3871 1266 3893
rect 1232 3825 1266 3833
rect 1232 3799 1266 3825
rect 1232 3757 1266 3761
rect 1232 3727 1266 3757
rect 1232 3655 1266 3689
rect 1232 3587 1266 3617
rect 1232 3583 1266 3587
rect 1232 3519 1266 3545
rect 1232 3511 1266 3519
rect 1232 3451 1266 3473
rect 1232 3439 1266 3451
rect 1232 3383 1266 3401
rect 1232 3367 1266 3383
rect 1232 3315 1266 3329
rect 1232 3295 1266 3315
rect 1232 3247 1266 3257
rect 1232 3223 1266 3247
rect 1232 3179 1266 3185
rect 1232 3151 1266 3179
rect 1232 3111 1266 3113
rect 1232 3079 1266 3111
rect 1232 3009 1266 3041
rect 1232 3007 1266 3009
rect 1232 2941 1266 2969
rect 1232 2935 1266 2941
rect 1232 2873 1266 2897
rect 1232 2863 1266 2873
rect 1232 2805 1266 2825
rect 1232 2791 1266 2805
rect 1232 2737 1266 2753
rect 1232 2719 1266 2737
rect 1232 2669 1266 2681
rect 1232 2647 1266 2669
rect 1232 2601 1266 2609
rect 1232 2575 1266 2601
rect 1232 2533 1266 2537
rect 1232 2503 1266 2533
rect 1232 2431 1266 2465
rect 1232 2363 1266 2393
rect 1232 2359 1266 2363
rect 1232 2295 1266 2321
rect 1232 2287 1266 2295
rect 1232 2227 1266 2249
rect 1232 2215 1266 2227
rect 1232 2159 1266 2177
rect 1232 2143 1266 2159
rect 1232 2091 1266 2105
rect 1232 2071 1266 2091
rect 1232 2023 1266 2033
rect 1232 1999 1266 2023
rect 1232 1955 1266 1961
rect 1232 1927 1266 1955
rect 1232 1887 1266 1889
rect 1232 1855 1266 1887
rect 1232 1785 1266 1817
rect 1232 1783 1266 1785
rect 1232 1717 1266 1745
rect 1232 1711 1266 1717
rect 1232 1649 1266 1673
rect 1232 1639 1266 1649
rect 1232 1581 1266 1601
rect 1232 1567 1266 1581
rect 1232 1513 1266 1529
rect 1232 1495 1266 1513
rect 1232 1445 1266 1457
rect 1232 1423 1266 1445
rect 1232 1377 1266 1385
rect 1232 1351 1266 1377
rect 1232 1309 1266 1313
rect 1232 1279 1266 1309
rect 1232 1207 1266 1241
rect 1232 1139 1266 1169
rect 1232 1135 1266 1139
rect 1232 1071 1266 1097
rect 1232 1063 1266 1071
rect 1232 1003 1266 1025
rect 1232 991 1266 1003
rect 1232 935 1266 953
rect 1232 919 1266 935
rect 1232 867 1266 881
rect 1232 847 1266 867
rect 1232 799 1266 809
rect 1232 775 1266 799
rect 1232 731 1266 737
rect 1232 703 1266 731
rect 1232 663 1266 665
rect 1232 631 1266 663
rect 1232 561 1266 593
rect 1232 559 1266 561
rect 1232 493 1266 521
rect 1232 487 1266 493
rect 1232 425 1266 449
rect 1232 415 1266 425
rect 1232 357 1266 377
rect 1232 343 1266 357
rect 1232 289 1266 305
rect 1232 271 1266 289
rect 1232 221 1266 233
rect 1232 199 1266 221
rect 1232 153 1266 161
rect 1232 127 1266 153
rect 1232 85 1266 89
rect 1232 55 1266 85
rect 1232 -17 1266 17
rect 1232 -85 1266 -55
rect 1232 -89 1266 -85
rect 1232 -153 1266 -127
rect 1232 -161 1266 -153
rect 1232 -221 1266 -199
rect 1232 -233 1266 -221
rect 1232 -289 1266 -271
rect 1232 -305 1266 -289
rect 1232 -357 1266 -343
rect 1232 -377 1266 -357
rect 1232 -425 1266 -415
rect 1232 -449 1266 -425
rect 1232 -493 1266 -487
rect 1232 -521 1266 -493
rect 1232 -561 1266 -559
rect 1232 -593 1266 -561
rect 1232 -663 1266 -631
rect 1232 -665 1266 -663
rect 1232 -731 1266 -703
rect 1232 -737 1266 -731
rect 1232 -799 1266 -775
rect 1232 -809 1266 -799
rect 1232 -867 1266 -847
rect 1232 -881 1266 -867
rect 1232 -935 1266 -919
rect 1232 -953 1266 -935
rect 1232 -1003 1266 -991
rect 1232 -1025 1266 -1003
rect 1232 -1071 1266 -1063
rect 1232 -1097 1266 -1071
rect 1232 -1139 1266 -1135
rect 1232 -1169 1266 -1139
rect 1232 -1241 1266 -1207
rect 1232 -1309 1266 -1279
rect 1232 -1313 1266 -1309
rect 1232 -1377 1266 -1351
rect 1232 -1385 1266 -1377
rect 1232 -1445 1266 -1423
rect 1232 -1457 1266 -1445
rect 1232 -1513 1266 -1495
rect 1232 -1529 1266 -1513
rect 1232 -1581 1266 -1567
rect 1232 -1601 1266 -1581
rect 1232 -1649 1266 -1639
rect 1232 -1673 1266 -1649
rect 1232 -1717 1266 -1711
rect 1232 -1745 1266 -1717
rect 1232 -1785 1266 -1783
rect 1232 -1817 1266 -1785
rect 1232 -1887 1266 -1855
rect 1232 -1889 1266 -1887
rect 1232 -1955 1266 -1927
rect 1232 -1961 1266 -1955
rect 1232 -2023 1266 -1999
rect 1232 -2033 1266 -2023
rect 1232 -2091 1266 -2071
rect 1232 -2105 1266 -2091
rect 1232 -2159 1266 -2143
rect 1232 -2177 1266 -2159
rect 1232 -2227 1266 -2215
rect 1232 -2249 1266 -2227
rect 1232 -2295 1266 -2287
rect 1232 -2321 1266 -2295
rect 1232 -2363 1266 -2359
rect 1232 -2393 1266 -2363
rect 1232 -2465 1266 -2431
rect 1232 -2533 1266 -2503
rect 1232 -2537 1266 -2533
rect 1232 -2601 1266 -2575
rect 1232 -2609 1266 -2601
rect 1232 -2669 1266 -2647
rect 1232 -2681 1266 -2669
rect 1232 -2737 1266 -2719
rect 1232 -2753 1266 -2737
rect 1232 -2805 1266 -2791
rect 1232 -2825 1266 -2805
rect 1232 -2873 1266 -2863
rect 1232 -2897 1266 -2873
rect 1232 -2941 1266 -2935
rect 1232 -2969 1266 -2941
rect 1232 -3009 1266 -3007
rect 1232 -3041 1266 -3009
rect 1232 -3111 1266 -3079
rect 1232 -3113 1266 -3111
rect 1232 -3179 1266 -3151
rect 1232 -3185 1266 -3179
rect 1232 -3247 1266 -3223
rect 1232 -3257 1266 -3247
rect 1232 -3315 1266 -3295
rect 1232 -3329 1266 -3315
rect 1232 -3383 1266 -3367
rect 1232 -3401 1266 -3383
rect 1232 -3451 1266 -3439
rect 1232 -3473 1266 -3451
rect 1232 -3519 1266 -3511
rect 1232 -3545 1266 -3519
rect 1232 -3587 1266 -3583
rect 1232 -3617 1266 -3587
rect 1232 -3689 1266 -3655
rect 1232 -3757 1266 -3727
rect 1232 -3761 1266 -3757
rect 1232 -3825 1266 -3799
rect 1232 -3833 1266 -3825
rect 1232 -3893 1266 -3871
rect 1232 -3905 1266 -3893
rect 1232 -3961 1266 -3943
rect 1232 -3977 1266 -3961
rect 1232 -4029 1266 -4015
rect 1232 -4049 1266 -4029
rect 1232 -4097 1266 -4087
rect 1232 -4121 1266 -4097
rect 1232 -4165 1266 -4159
rect 1232 -4193 1266 -4165
rect 1232 -4233 1266 -4231
rect 1232 -4265 1266 -4233
rect 1232 -4335 1266 -4303
rect 1232 -4337 1266 -4335
rect 1232 -4403 1266 -4375
rect 1232 -4409 1266 -4403
rect 1232 -4471 1266 -4447
rect 1232 -4481 1266 -4471
rect 1232 -4539 1266 -4519
rect 1232 -4553 1266 -4539
rect 1232 -4607 1266 -4591
rect 1232 -4625 1266 -4607
rect 1232 -4675 1266 -4663
rect 1232 -4697 1266 -4675
rect 1232 -4743 1266 -4735
rect 1232 -4769 1266 -4743
rect 1232 -4811 1266 -4807
rect 1232 -4841 1266 -4811
rect 1232 -4913 1266 -4879
rect 1232 -4981 1266 -4951
rect 1232 -4985 1266 -4981
rect -1153 -5102 -1149 -5068
rect -1149 -5102 -1119 -5068
rect -1081 -5102 -1047 -5068
rect -1009 -5102 -979 -5068
rect -979 -5102 -975 -5068
rect -621 -5102 -617 -5068
rect -617 -5102 -587 -5068
rect -549 -5102 -515 -5068
rect -477 -5102 -447 -5068
rect -447 -5102 -443 -5068
rect -89 -5102 -85 -5068
rect -85 -5102 -55 -5068
rect -17 -5102 17 -5068
rect 55 -5102 85 -5068
rect 85 -5102 89 -5068
rect 443 -5102 447 -5068
rect 447 -5102 477 -5068
rect 515 -5102 549 -5068
rect 587 -5102 617 -5068
rect 617 -5102 621 -5068
rect 975 -5102 979 -5068
rect 979 -5102 1009 -5068
rect 1047 -5102 1081 -5068
rect 1119 -5102 1149 -5068
rect 1149 -5102 1153 -5068
rect 1542 5219 1936 5237
rect 1542 -5219 1552 5219
rect 1552 -5219 1926 5219
rect 1926 -5219 1936 5219
rect 1542 -5237 1936 -5219
rect -1421 -5356 1421 -5346
rect -1421 -5730 -1411 -5356
rect -1411 -5730 1411 -5356
rect 1411 -5730 1421 -5356
rect -1421 -5740 1421 -5730
<< metal1 >>
tri -1576 5740 -1556 5760 se
rect -1556 5740 1556 5760
tri -1956 5360 -1576 5740 se
rect -1576 5360 -1421 5740
rect -1956 5346 -1421 5360
rect 1421 5360 1556 5740
tri 1556 5360 1956 5760 sw
rect 1421 5346 1956 5360
rect -1956 5295 1956 5346
rect -1956 5268 -1480 5295
tri -1480 5268 -1453 5295 nw
tri 1448 5268 1475 5295 ne
rect 1475 5268 1956 5295
rect -1956 5237 -1493 5268
tri -1493 5255 -1480 5268 nw
tri 1475 5255 1488 5268 ne
rect -1956 -5237 -1936 5237
rect -1542 -5237 -1493 5237
rect 1488 5237 1956 5268
rect -1330 5102 1330 5168
rect -1330 5068 -1153 5102
rect -1119 5068 -1081 5102
rect -1047 5068 -1009 5102
rect -975 5068 -621 5102
rect -587 5068 -549 5102
rect -515 5068 -477 5102
rect -443 5068 -89 5102
rect -55 5068 -17 5102
rect 17 5068 55 5102
rect 89 5068 443 5102
rect 477 5068 515 5102
rect 549 5068 587 5102
rect 621 5068 975 5102
rect 1009 5068 1047 5102
rect 1081 5068 1119 5102
rect 1153 5068 1330 5102
rect -1330 5062 1330 5068
rect -1330 4985 -1226 5062
tri -1226 5022 -1186 5062 nw
tri -942 5022 -902 5062 ne
rect -1330 4951 -1266 4985
rect -1232 4951 -1226 4985
rect -1330 4913 -1226 4951
rect -1330 4879 -1266 4913
rect -1232 4879 -1226 4913
rect -1330 4841 -1226 4879
rect -1330 4807 -1266 4841
rect -1232 4807 -1226 4841
rect -1330 4769 -1226 4807
rect -1330 4735 -1266 4769
rect -1232 4735 -1226 4769
rect -1330 4697 -1226 4735
rect -1330 4663 -1266 4697
rect -1232 4663 -1226 4697
rect -1330 4625 -1226 4663
rect -1330 4591 -1266 4625
rect -1232 4591 -1226 4625
rect -1330 4553 -1226 4591
rect -1330 4519 -1266 4553
rect -1232 4519 -1226 4553
rect -1330 4481 -1226 4519
rect -1330 4447 -1266 4481
rect -1232 4447 -1226 4481
rect -1330 4409 -1226 4447
rect -1330 4375 -1266 4409
rect -1232 4375 -1226 4409
rect -1330 4337 -1226 4375
rect -1330 4303 -1266 4337
rect -1232 4303 -1226 4337
rect -1330 4265 -1226 4303
rect -1330 4231 -1266 4265
rect -1232 4231 -1226 4265
rect -1330 4193 -1226 4231
rect -1330 4159 -1266 4193
rect -1232 4159 -1226 4193
rect -1330 4121 -1226 4159
rect -1330 4087 -1266 4121
rect -1232 4087 -1226 4121
rect -1330 4049 -1226 4087
rect -1330 4015 -1266 4049
rect -1232 4015 -1226 4049
rect -1330 3977 -1226 4015
rect -1330 3943 -1266 3977
rect -1232 3943 -1226 3977
rect -1330 3905 -1226 3943
rect -1330 3871 -1266 3905
rect -1232 3871 -1226 3905
rect -1330 3833 -1226 3871
rect -1330 3799 -1266 3833
rect -1232 3799 -1226 3833
rect -1330 3761 -1226 3799
rect -1330 3727 -1266 3761
rect -1232 3727 -1226 3761
rect -1330 3689 -1226 3727
rect -1330 3655 -1266 3689
rect -1232 3655 -1226 3689
rect -1330 3617 -1226 3655
rect -1330 3583 -1266 3617
rect -1232 3583 -1226 3617
rect -1330 3545 -1226 3583
rect -1330 3511 -1266 3545
rect -1232 3511 -1226 3545
rect -1330 3473 -1226 3511
rect -1330 3439 -1266 3473
rect -1232 3439 -1226 3473
rect -1330 3401 -1226 3439
rect -1330 3367 -1266 3401
rect -1232 3367 -1226 3401
rect -1330 3329 -1226 3367
rect -1330 3295 -1266 3329
rect -1232 3295 -1226 3329
rect -1330 3257 -1226 3295
rect -1330 3223 -1266 3257
rect -1232 3223 -1226 3257
rect -1330 3185 -1226 3223
rect -1330 3151 -1266 3185
rect -1232 3151 -1226 3185
rect -1330 3113 -1226 3151
rect -1330 3079 -1266 3113
rect -1232 3079 -1226 3113
rect -1330 3041 -1226 3079
rect -1330 3007 -1266 3041
rect -1232 3007 -1226 3041
rect -1330 2969 -1226 3007
rect -1330 2935 -1266 2969
rect -1232 2935 -1226 2969
rect -1330 2897 -1226 2935
rect -1330 2863 -1266 2897
rect -1232 2863 -1226 2897
rect -1330 2825 -1226 2863
rect -1330 2791 -1266 2825
rect -1232 2791 -1226 2825
rect -1330 2753 -1226 2791
rect -1330 2719 -1266 2753
rect -1232 2719 -1226 2753
rect -1330 2681 -1226 2719
rect -1330 2647 -1266 2681
rect -1232 2647 -1226 2681
rect -1330 2609 -1226 2647
rect -1330 2575 -1266 2609
rect -1232 2575 -1226 2609
rect -1330 2537 -1226 2575
rect -1330 2503 -1266 2537
rect -1232 2503 -1226 2537
rect -1330 2465 -1226 2503
rect -1330 2431 -1266 2465
rect -1232 2431 -1226 2465
rect -1330 2393 -1226 2431
rect -1330 2359 -1266 2393
rect -1232 2359 -1226 2393
rect -1330 2321 -1226 2359
rect -1330 2287 -1266 2321
rect -1232 2287 -1226 2321
rect -1330 2249 -1226 2287
rect -1330 2215 -1266 2249
rect -1232 2215 -1226 2249
rect -1330 2177 -1226 2215
rect -1330 2143 -1266 2177
rect -1232 2143 -1226 2177
rect -1330 2105 -1226 2143
rect -1330 2071 -1266 2105
rect -1232 2071 -1226 2105
rect -1330 2033 -1226 2071
rect -1330 1999 -1266 2033
rect -1232 1999 -1226 2033
rect -1330 1961 -1226 1999
rect -1330 1927 -1266 1961
rect -1232 1927 -1226 1961
rect -1330 1889 -1226 1927
rect -1330 1855 -1266 1889
rect -1232 1855 -1226 1889
rect -1330 1817 -1226 1855
rect -1330 1783 -1266 1817
rect -1232 1783 -1226 1817
rect -1330 1745 -1226 1783
rect -1330 1711 -1266 1745
rect -1232 1711 -1226 1745
rect -1330 1673 -1226 1711
rect -1330 1639 -1266 1673
rect -1232 1639 -1226 1673
rect -1330 1601 -1226 1639
rect -1330 1567 -1266 1601
rect -1232 1567 -1226 1601
rect -1330 1529 -1226 1567
rect -1330 1495 -1266 1529
rect -1232 1495 -1226 1529
rect -1330 1457 -1226 1495
rect -1330 1423 -1266 1457
rect -1232 1423 -1226 1457
rect -1330 1385 -1226 1423
rect -1330 1351 -1266 1385
rect -1232 1351 -1226 1385
rect -1330 1313 -1226 1351
rect -1330 1279 -1266 1313
rect -1232 1279 -1226 1313
rect -1330 1241 -1226 1279
rect -1330 1207 -1266 1241
rect -1232 1207 -1226 1241
rect -1330 1169 -1226 1207
rect -1330 1135 -1266 1169
rect -1232 1135 -1226 1169
rect -1330 1097 -1226 1135
rect -1330 1063 -1266 1097
rect -1232 1063 -1226 1097
rect -1330 1025 -1226 1063
rect -1330 991 -1266 1025
rect -1232 991 -1226 1025
rect -1330 953 -1226 991
rect -1330 919 -1266 953
rect -1232 919 -1226 953
rect -1330 881 -1226 919
rect -1330 847 -1266 881
rect -1232 847 -1226 881
rect -1330 809 -1226 847
rect -1330 775 -1266 809
rect -1232 775 -1226 809
rect -1330 737 -1226 775
rect -1330 703 -1266 737
rect -1232 703 -1226 737
rect -1330 665 -1226 703
rect -1330 631 -1266 665
rect -1232 631 -1226 665
rect -1330 593 -1226 631
rect -1330 559 -1266 593
rect -1232 559 -1226 593
rect -1330 521 -1226 559
rect -1330 487 -1266 521
rect -1232 487 -1226 521
rect -1330 449 -1226 487
rect -1330 415 -1266 449
rect -1232 415 -1226 449
rect -1330 377 -1226 415
rect -1330 343 -1266 377
rect -1232 343 -1226 377
rect -1330 305 -1226 343
rect -1330 271 -1266 305
rect -1232 271 -1226 305
rect -1330 233 -1226 271
rect -1330 199 -1266 233
rect -1232 199 -1226 233
rect -1330 161 -1226 199
rect -1330 127 -1266 161
rect -1232 127 -1226 161
rect -1330 89 -1226 127
rect -1330 55 -1266 89
rect -1232 55 -1226 89
rect -1330 17 -1226 55
rect -1330 -17 -1266 17
rect -1232 -17 -1226 17
rect -1330 -55 -1226 -17
rect -1330 -89 -1266 -55
rect -1232 -89 -1226 -55
rect -1330 -127 -1226 -89
rect -1330 -161 -1266 -127
rect -1232 -161 -1226 -127
rect -1330 -199 -1226 -161
rect -1330 -233 -1266 -199
rect -1232 -233 -1226 -199
rect -1330 -271 -1226 -233
rect -1330 -305 -1266 -271
rect -1232 -305 -1226 -271
rect -1330 -343 -1226 -305
rect -1330 -377 -1266 -343
rect -1232 -377 -1226 -343
rect -1330 -415 -1226 -377
rect -1330 -449 -1266 -415
rect -1232 -449 -1226 -415
rect -1330 -487 -1226 -449
rect -1330 -521 -1266 -487
rect -1232 -521 -1226 -487
rect -1330 -559 -1226 -521
rect -1330 -593 -1266 -559
rect -1232 -593 -1226 -559
rect -1330 -631 -1226 -593
rect -1330 -665 -1266 -631
rect -1232 -665 -1226 -631
rect -1330 -703 -1226 -665
rect -1330 -737 -1266 -703
rect -1232 -737 -1226 -703
rect -1330 -775 -1226 -737
rect -1330 -809 -1266 -775
rect -1232 -809 -1226 -775
rect -1330 -847 -1226 -809
rect -1330 -881 -1266 -847
rect -1232 -881 -1226 -847
rect -1330 -919 -1226 -881
rect -1330 -953 -1266 -919
rect -1232 -953 -1226 -919
rect -1330 -991 -1226 -953
rect -1330 -1025 -1266 -991
rect -1232 -1025 -1226 -991
rect -1330 -1063 -1226 -1025
rect -1330 -1097 -1266 -1063
rect -1232 -1097 -1226 -1063
rect -1330 -1135 -1226 -1097
rect -1330 -1169 -1266 -1135
rect -1232 -1169 -1226 -1135
rect -1330 -1207 -1226 -1169
rect -1330 -1241 -1266 -1207
rect -1232 -1241 -1226 -1207
rect -1330 -1279 -1226 -1241
rect -1330 -1313 -1266 -1279
rect -1232 -1313 -1226 -1279
rect -1330 -1351 -1226 -1313
rect -1330 -1385 -1266 -1351
rect -1232 -1385 -1226 -1351
rect -1330 -1423 -1226 -1385
rect -1330 -1457 -1266 -1423
rect -1232 -1457 -1226 -1423
rect -1330 -1495 -1226 -1457
rect -1330 -1529 -1266 -1495
rect -1232 -1529 -1226 -1495
rect -1330 -1567 -1226 -1529
rect -1330 -1601 -1266 -1567
rect -1232 -1601 -1226 -1567
rect -1330 -1639 -1226 -1601
rect -1330 -1673 -1266 -1639
rect -1232 -1673 -1226 -1639
rect -1330 -1711 -1226 -1673
rect -1330 -1745 -1266 -1711
rect -1232 -1745 -1226 -1711
rect -1330 -1783 -1226 -1745
rect -1330 -1817 -1266 -1783
rect -1232 -1817 -1226 -1783
rect -1330 -1855 -1226 -1817
rect -1330 -1889 -1266 -1855
rect -1232 -1889 -1226 -1855
rect -1330 -1927 -1226 -1889
rect -1330 -1961 -1266 -1927
rect -1232 -1961 -1226 -1927
rect -1330 -1999 -1226 -1961
rect -1330 -2033 -1266 -1999
rect -1232 -2033 -1226 -1999
rect -1330 -2071 -1226 -2033
rect -1330 -2105 -1266 -2071
rect -1232 -2105 -1226 -2071
rect -1330 -2143 -1226 -2105
rect -1330 -2177 -1266 -2143
rect -1232 -2177 -1226 -2143
rect -1330 -2215 -1226 -2177
rect -1330 -2249 -1266 -2215
rect -1232 -2249 -1226 -2215
rect -1330 -2287 -1226 -2249
rect -1330 -2321 -1266 -2287
rect -1232 -2321 -1226 -2287
rect -1330 -2359 -1226 -2321
rect -1330 -2393 -1266 -2359
rect -1232 -2393 -1226 -2359
rect -1330 -2431 -1226 -2393
rect -1330 -2465 -1266 -2431
rect -1232 -2465 -1226 -2431
rect -1330 -2503 -1226 -2465
rect -1330 -2537 -1266 -2503
rect -1232 -2537 -1226 -2503
rect -1330 -2575 -1226 -2537
rect -1330 -2609 -1266 -2575
rect -1232 -2609 -1226 -2575
rect -1330 -2647 -1226 -2609
rect -1330 -2681 -1266 -2647
rect -1232 -2681 -1226 -2647
rect -1330 -2719 -1226 -2681
rect -1330 -2753 -1266 -2719
rect -1232 -2753 -1226 -2719
rect -1330 -2791 -1226 -2753
rect -1330 -2825 -1266 -2791
rect -1232 -2825 -1226 -2791
rect -1330 -2863 -1226 -2825
rect -1330 -2897 -1266 -2863
rect -1232 -2897 -1226 -2863
rect -1330 -2935 -1226 -2897
rect -1330 -2969 -1266 -2935
rect -1232 -2969 -1226 -2935
rect -1330 -3007 -1226 -2969
rect -1330 -3041 -1266 -3007
rect -1232 -3041 -1226 -3007
rect -1330 -3079 -1226 -3041
rect -1330 -3113 -1266 -3079
rect -1232 -3113 -1226 -3079
rect -1330 -3151 -1226 -3113
rect -1330 -3185 -1266 -3151
rect -1232 -3185 -1226 -3151
rect -1330 -3223 -1226 -3185
rect -1330 -3257 -1266 -3223
rect -1232 -3257 -1226 -3223
rect -1330 -3295 -1226 -3257
rect -1330 -3329 -1266 -3295
rect -1232 -3329 -1226 -3295
rect -1330 -3367 -1226 -3329
rect -1330 -3401 -1266 -3367
rect -1232 -3401 -1226 -3367
rect -1330 -3439 -1226 -3401
rect -1330 -3473 -1266 -3439
rect -1232 -3473 -1226 -3439
rect -1330 -3511 -1226 -3473
rect -1330 -3545 -1266 -3511
rect -1232 -3545 -1226 -3511
rect -1330 -3583 -1226 -3545
rect -1330 -3617 -1266 -3583
rect -1232 -3617 -1226 -3583
rect -1330 -3655 -1226 -3617
rect -1330 -3689 -1266 -3655
rect -1232 -3689 -1226 -3655
rect -1330 -3727 -1226 -3689
rect -1330 -3761 -1266 -3727
rect -1232 -3761 -1226 -3727
rect -1330 -3799 -1226 -3761
rect -1330 -3833 -1266 -3799
rect -1232 -3833 -1226 -3799
rect -1330 -3871 -1226 -3833
rect -1330 -3905 -1266 -3871
rect -1232 -3905 -1226 -3871
rect -1330 -3943 -1226 -3905
rect -1330 -3977 -1266 -3943
rect -1232 -3977 -1226 -3943
rect -1330 -4015 -1226 -3977
rect -1330 -4049 -1266 -4015
rect -1232 -4049 -1226 -4015
rect -1330 -4087 -1226 -4049
rect -1330 -4121 -1266 -4087
rect -1232 -4121 -1226 -4087
rect -1330 -4159 -1226 -4121
rect -1330 -4193 -1266 -4159
rect -1232 -4193 -1226 -4159
rect -1330 -4231 -1226 -4193
rect -1330 -4265 -1266 -4231
rect -1232 -4265 -1226 -4231
rect -1330 -4303 -1226 -4265
rect -1330 -4337 -1266 -4303
rect -1232 -4337 -1226 -4303
rect -1330 -4375 -1226 -4337
rect -1330 -4409 -1266 -4375
rect -1232 -4409 -1226 -4375
rect -1330 -4447 -1226 -4409
rect -1330 -4481 -1266 -4447
rect -1232 -4481 -1226 -4447
rect -1330 -4519 -1226 -4481
rect -1330 -4553 -1266 -4519
rect -1232 -4553 -1226 -4519
rect -1330 -4591 -1226 -4553
rect -1330 -4625 -1266 -4591
rect -1232 -4625 -1226 -4591
rect -1330 -4663 -1226 -4625
rect -1330 -4697 -1266 -4663
rect -1232 -4697 -1226 -4663
rect -1330 -4735 -1226 -4697
rect -1330 -4769 -1266 -4735
rect -1232 -4769 -1226 -4735
rect -1330 -4807 -1226 -4769
rect -1330 -4841 -1266 -4807
rect -1232 -4841 -1226 -4807
rect -1330 -4879 -1226 -4841
rect -1330 -4913 -1266 -4879
rect -1232 -4913 -1226 -4879
rect -1330 -4951 -1226 -4913
rect -1330 -4985 -1266 -4951
rect -1232 -4985 -1226 -4951
rect -1330 -5062 -1226 -4985
tri -1158 5000 -1138 5020 se
rect -1138 5000 -990 5020
tri -990 5000 -970 5020 sw
rect -1158 4985 -970 5000
rect -1158 -4985 -1117 4985
rect -1011 -4985 -970 4985
rect -1158 -5000 -970 -4985
tri -1158 -5020 -1138 -5000 ne
rect -1138 -5020 -990 -5000
tri -990 -5020 -970 -5000 nw
rect -902 4985 -694 5062
tri -694 5022 -654 5062 nw
tri -410 5022 -370 5062 ne
rect -902 4951 -896 4985
rect -862 4951 -815 4985
rect -781 4951 -734 4985
rect -700 4951 -694 4985
rect -902 4913 -694 4951
rect -902 4879 -896 4913
rect -862 4879 -815 4913
rect -781 4879 -734 4913
rect -700 4879 -694 4913
rect -902 4841 -694 4879
rect -902 4807 -896 4841
rect -862 4807 -815 4841
rect -781 4807 -734 4841
rect -700 4807 -694 4841
rect -902 4769 -694 4807
rect -902 4735 -896 4769
rect -862 4735 -815 4769
rect -781 4735 -734 4769
rect -700 4735 -694 4769
rect -902 4697 -694 4735
rect -902 4663 -896 4697
rect -862 4663 -815 4697
rect -781 4663 -734 4697
rect -700 4663 -694 4697
rect -902 4625 -694 4663
rect -902 4591 -896 4625
rect -862 4591 -815 4625
rect -781 4591 -734 4625
rect -700 4591 -694 4625
rect -902 4553 -694 4591
rect -902 4519 -896 4553
rect -862 4519 -815 4553
rect -781 4519 -734 4553
rect -700 4519 -694 4553
rect -902 4481 -694 4519
rect -902 4447 -896 4481
rect -862 4447 -815 4481
rect -781 4447 -734 4481
rect -700 4447 -694 4481
rect -902 4409 -694 4447
rect -902 4375 -896 4409
rect -862 4375 -815 4409
rect -781 4375 -734 4409
rect -700 4375 -694 4409
rect -902 4337 -694 4375
rect -902 4303 -896 4337
rect -862 4303 -815 4337
rect -781 4303 -734 4337
rect -700 4303 -694 4337
rect -902 4265 -694 4303
rect -902 4231 -896 4265
rect -862 4231 -815 4265
rect -781 4231 -734 4265
rect -700 4231 -694 4265
rect -902 4193 -694 4231
rect -902 4159 -896 4193
rect -862 4159 -815 4193
rect -781 4159 -734 4193
rect -700 4159 -694 4193
rect -902 4121 -694 4159
rect -902 4087 -896 4121
rect -862 4087 -815 4121
rect -781 4087 -734 4121
rect -700 4087 -694 4121
rect -902 4049 -694 4087
rect -902 4015 -896 4049
rect -862 4015 -815 4049
rect -781 4015 -734 4049
rect -700 4015 -694 4049
rect -902 3977 -694 4015
rect -902 3943 -896 3977
rect -862 3943 -815 3977
rect -781 3943 -734 3977
rect -700 3943 -694 3977
rect -902 3905 -694 3943
rect -902 3871 -896 3905
rect -862 3871 -815 3905
rect -781 3871 -734 3905
rect -700 3871 -694 3905
rect -902 3833 -694 3871
rect -902 3799 -896 3833
rect -862 3799 -815 3833
rect -781 3799 -734 3833
rect -700 3799 -694 3833
rect -902 3761 -694 3799
rect -902 3727 -896 3761
rect -862 3727 -815 3761
rect -781 3727 -734 3761
rect -700 3727 -694 3761
rect -902 3689 -694 3727
rect -902 3655 -896 3689
rect -862 3655 -815 3689
rect -781 3655 -734 3689
rect -700 3655 -694 3689
rect -902 3617 -694 3655
rect -902 3583 -896 3617
rect -862 3583 -815 3617
rect -781 3583 -734 3617
rect -700 3583 -694 3617
rect -902 3545 -694 3583
rect -902 3511 -896 3545
rect -862 3511 -815 3545
rect -781 3511 -734 3545
rect -700 3511 -694 3545
rect -902 3473 -694 3511
rect -902 3439 -896 3473
rect -862 3439 -815 3473
rect -781 3439 -734 3473
rect -700 3439 -694 3473
rect -902 3401 -694 3439
rect -902 3367 -896 3401
rect -862 3367 -815 3401
rect -781 3367 -734 3401
rect -700 3367 -694 3401
rect -902 3329 -694 3367
rect -902 3295 -896 3329
rect -862 3295 -815 3329
rect -781 3295 -734 3329
rect -700 3295 -694 3329
rect -902 3257 -694 3295
rect -902 3223 -896 3257
rect -862 3223 -815 3257
rect -781 3223 -734 3257
rect -700 3223 -694 3257
rect -902 3185 -694 3223
rect -902 3151 -896 3185
rect -862 3151 -815 3185
rect -781 3151 -734 3185
rect -700 3151 -694 3185
rect -902 3113 -694 3151
rect -902 3079 -896 3113
rect -862 3079 -815 3113
rect -781 3079 -734 3113
rect -700 3079 -694 3113
rect -902 3041 -694 3079
rect -902 3007 -896 3041
rect -862 3007 -815 3041
rect -781 3007 -734 3041
rect -700 3007 -694 3041
rect -902 2969 -694 3007
rect -902 2935 -896 2969
rect -862 2935 -815 2969
rect -781 2935 -734 2969
rect -700 2935 -694 2969
rect -902 2897 -694 2935
rect -902 2863 -896 2897
rect -862 2863 -815 2897
rect -781 2863 -734 2897
rect -700 2863 -694 2897
rect -902 2825 -694 2863
rect -902 2791 -896 2825
rect -862 2791 -815 2825
rect -781 2791 -734 2825
rect -700 2791 -694 2825
rect -902 2753 -694 2791
rect -902 2719 -896 2753
rect -862 2719 -815 2753
rect -781 2719 -734 2753
rect -700 2719 -694 2753
rect -902 2681 -694 2719
rect -902 2647 -896 2681
rect -862 2647 -815 2681
rect -781 2647 -734 2681
rect -700 2647 -694 2681
rect -902 2609 -694 2647
rect -902 2575 -896 2609
rect -862 2575 -815 2609
rect -781 2575 -734 2609
rect -700 2575 -694 2609
rect -902 2537 -694 2575
rect -902 2503 -896 2537
rect -862 2503 -815 2537
rect -781 2503 -734 2537
rect -700 2503 -694 2537
rect -902 2465 -694 2503
rect -902 2431 -896 2465
rect -862 2431 -815 2465
rect -781 2431 -734 2465
rect -700 2431 -694 2465
rect -902 2393 -694 2431
rect -902 2359 -896 2393
rect -862 2359 -815 2393
rect -781 2359 -734 2393
rect -700 2359 -694 2393
rect -902 2321 -694 2359
rect -902 2287 -896 2321
rect -862 2287 -815 2321
rect -781 2287 -734 2321
rect -700 2287 -694 2321
rect -902 2249 -694 2287
rect -902 2215 -896 2249
rect -862 2215 -815 2249
rect -781 2215 -734 2249
rect -700 2215 -694 2249
rect -902 2177 -694 2215
rect -902 2143 -896 2177
rect -862 2143 -815 2177
rect -781 2143 -734 2177
rect -700 2143 -694 2177
rect -902 2105 -694 2143
rect -902 2071 -896 2105
rect -862 2071 -815 2105
rect -781 2071 -734 2105
rect -700 2071 -694 2105
rect -902 2033 -694 2071
rect -902 1999 -896 2033
rect -862 1999 -815 2033
rect -781 1999 -734 2033
rect -700 1999 -694 2033
rect -902 1961 -694 1999
rect -902 1927 -896 1961
rect -862 1927 -815 1961
rect -781 1927 -734 1961
rect -700 1927 -694 1961
rect -902 1889 -694 1927
rect -902 1855 -896 1889
rect -862 1855 -815 1889
rect -781 1855 -734 1889
rect -700 1855 -694 1889
rect -902 1817 -694 1855
rect -902 1783 -896 1817
rect -862 1783 -815 1817
rect -781 1783 -734 1817
rect -700 1783 -694 1817
rect -902 1745 -694 1783
rect -902 1711 -896 1745
rect -862 1711 -815 1745
rect -781 1711 -734 1745
rect -700 1711 -694 1745
rect -902 1673 -694 1711
rect -902 1639 -896 1673
rect -862 1639 -815 1673
rect -781 1639 -734 1673
rect -700 1639 -694 1673
rect -902 1601 -694 1639
rect -902 1567 -896 1601
rect -862 1567 -815 1601
rect -781 1567 -734 1601
rect -700 1567 -694 1601
rect -902 1529 -694 1567
rect -902 1495 -896 1529
rect -862 1495 -815 1529
rect -781 1495 -734 1529
rect -700 1495 -694 1529
rect -902 1457 -694 1495
rect -902 1423 -896 1457
rect -862 1423 -815 1457
rect -781 1423 -734 1457
rect -700 1423 -694 1457
rect -902 1385 -694 1423
rect -902 1351 -896 1385
rect -862 1351 -815 1385
rect -781 1351 -734 1385
rect -700 1351 -694 1385
rect -902 1313 -694 1351
rect -902 1279 -896 1313
rect -862 1279 -815 1313
rect -781 1279 -734 1313
rect -700 1279 -694 1313
rect -902 1241 -694 1279
rect -902 1207 -896 1241
rect -862 1207 -815 1241
rect -781 1207 -734 1241
rect -700 1207 -694 1241
rect -902 1169 -694 1207
rect -902 1135 -896 1169
rect -862 1135 -815 1169
rect -781 1135 -734 1169
rect -700 1135 -694 1169
rect -902 1097 -694 1135
rect -902 1063 -896 1097
rect -862 1063 -815 1097
rect -781 1063 -734 1097
rect -700 1063 -694 1097
rect -902 1025 -694 1063
rect -902 991 -896 1025
rect -862 991 -815 1025
rect -781 991 -734 1025
rect -700 991 -694 1025
rect -902 953 -694 991
rect -902 919 -896 953
rect -862 919 -815 953
rect -781 919 -734 953
rect -700 919 -694 953
rect -902 881 -694 919
rect -902 847 -896 881
rect -862 847 -815 881
rect -781 847 -734 881
rect -700 847 -694 881
rect -902 809 -694 847
rect -902 775 -896 809
rect -862 775 -815 809
rect -781 775 -734 809
rect -700 775 -694 809
rect -902 737 -694 775
rect -902 703 -896 737
rect -862 703 -815 737
rect -781 703 -734 737
rect -700 703 -694 737
rect -902 665 -694 703
rect -902 631 -896 665
rect -862 631 -815 665
rect -781 631 -734 665
rect -700 631 -694 665
rect -902 593 -694 631
rect -902 559 -896 593
rect -862 559 -815 593
rect -781 559 -734 593
rect -700 559 -694 593
rect -902 521 -694 559
rect -902 487 -896 521
rect -862 487 -815 521
rect -781 487 -734 521
rect -700 487 -694 521
rect -902 449 -694 487
rect -902 415 -896 449
rect -862 415 -815 449
rect -781 415 -734 449
rect -700 415 -694 449
rect -902 377 -694 415
rect -902 343 -896 377
rect -862 343 -815 377
rect -781 343 -734 377
rect -700 343 -694 377
rect -902 305 -694 343
rect -902 271 -896 305
rect -862 271 -815 305
rect -781 271 -734 305
rect -700 271 -694 305
rect -902 233 -694 271
rect -902 199 -896 233
rect -862 199 -815 233
rect -781 199 -734 233
rect -700 199 -694 233
rect -902 161 -694 199
rect -902 127 -896 161
rect -862 127 -815 161
rect -781 127 -734 161
rect -700 127 -694 161
rect -902 89 -694 127
rect -902 55 -896 89
rect -862 55 -815 89
rect -781 55 -734 89
rect -700 55 -694 89
rect -902 17 -694 55
rect -902 -17 -896 17
rect -862 -17 -815 17
rect -781 -17 -734 17
rect -700 -17 -694 17
rect -902 -55 -694 -17
rect -902 -89 -896 -55
rect -862 -89 -815 -55
rect -781 -89 -734 -55
rect -700 -89 -694 -55
rect -902 -127 -694 -89
rect -902 -161 -896 -127
rect -862 -161 -815 -127
rect -781 -161 -734 -127
rect -700 -161 -694 -127
rect -902 -199 -694 -161
rect -902 -233 -896 -199
rect -862 -233 -815 -199
rect -781 -233 -734 -199
rect -700 -233 -694 -199
rect -902 -271 -694 -233
rect -902 -305 -896 -271
rect -862 -305 -815 -271
rect -781 -305 -734 -271
rect -700 -305 -694 -271
rect -902 -343 -694 -305
rect -902 -377 -896 -343
rect -862 -377 -815 -343
rect -781 -377 -734 -343
rect -700 -377 -694 -343
rect -902 -415 -694 -377
rect -902 -449 -896 -415
rect -862 -449 -815 -415
rect -781 -449 -734 -415
rect -700 -449 -694 -415
rect -902 -487 -694 -449
rect -902 -521 -896 -487
rect -862 -521 -815 -487
rect -781 -521 -734 -487
rect -700 -521 -694 -487
rect -902 -559 -694 -521
rect -902 -593 -896 -559
rect -862 -593 -815 -559
rect -781 -593 -734 -559
rect -700 -593 -694 -559
rect -902 -631 -694 -593
rect -902 -665 -896 -631
rect -862 -665 -815 -631
rect -781 -665 -734 -631
rect -700 -665 -694 -631
rect -902 -703 -694 -665
rect -902 -737 -896 -703
rect -862 -737 -815 -703
rect -781 -737 -734 -703
rect -700 -737 -694 -703
rect -902 -775 -694 -737
rect -902 -809 -896 -775
rect -862 -809 -815 -775
rect -781 -809 -734 -775
rect -700 -809 -694 -775
rect -902 -847 -694 -809
rect -902 -881 -896 -847
rect -862 -881 -815 -847
rect -781 -881 -734 -847
rect -700 -881 -694 -847
rect -902 -919 -694 -881
rect -902 -953 -896 -919
rect -862 -953 -815 -919
rect -781 -953 -734 -919
rect -700 -953 -694 -919
rect -902 -991 -694 -953
rect -902 -1025 -896 -991
rect -862 -1025 -815 -991
rect -781 -1025 -734 -991
rect -700 -1025 -694 -991
rect -902 -1063 -694 -1025
rect -902 -1097 -896 -1063
rect -862 -1097 -815 -1063
rect -781 -1097 -734 -1063
rect -700 -1097 -694 -1063
rect -902 -1135 -694 -1097
rect -902 -1169 -896 -1135
rect -862 -1169 -815 -1135
rect -781 -1169 -734 -1135
rect -700 -1169 -694 -1135
rect -902 -1207 -694 -1169
rect -902 -1241 -896 -1207
rect -862 -1241 -815 -1207
rect -781 -1241 -734 -1207
rect -700 -1241 -694 -1207
rect -902 -1279 -694 -1241
rect -902 -1313 -896 -1279
rect -862 -1313 -815 -1279
rect -781 -1313 -734 -1279
rect -700 -1313 -694 -1279
rect -902 -1351 -694 -1313
rect -902 -1385 -896 -1351
rect -862 -1385 -815 -1351
rect -781 -1385 -734 -1351
rect -700 -1385 -694 -1351
rect -902 -1423 -694 -1385
rect -902 -1457 -896 -1423
rect -862 -1457 -815 -1423
rect -781 -1457 -734 -1423
rect -700 -1457 -694 -1423
rect -902 -1495 -694 -1457
rect -902 -1529 -896 -1495
rect -862 -1529 -815 -1495
rect -781 -1529 -734 -1495
rect -700 -1529 -694 -1495
rect -902 -1567 -694 -1529
rect -902 -1601 -896 -1567
rect -862 -1601 -815 -1567
rect -781 -1601 -734 -1567
rect -700 -1601 -694 -1567
rect -902 -1639 -694 -1601
rect -902 -1673 -896 -1639
rect -862 -1673 -815 -1639
rect -781 -1673 -734 -1639
rect -700 -1673 -694 -1639
rect -902 -1711 -694 -1673
rect -902 -1745 -896 -1711
rect -862 -1745 -815 -1711
rect -781 -1745 -734 -1711
rect -700 -1745 -694 -1711
rect -902 -1783 -694 -1745
rect -902 -1817 -896 -1783
rect -862 -1817 -815 -1783
rect -781 -1817 -734 -1783
rect -700 -1817 -694 -1783
rect -902 -1855 -694 -1817
rect -902 -1889 -896 -1855
rect -862 -1889 -815 -1855
rect -781 -1889 -734 -1855
rect -700 -1889 -694 -1855
rect -902 -1927 -694 -1889
rect -902 -1961 -896 -1927
rect -862 -1961 -815 -1927
rect -781 -1961 -734 -1927
rect -700 -1961 -694 -1927
rect -902 -1999 -694 -1961
rect -902 -2033 -896 -1999
rect -862 -2033 -815 -1999
rect -781 -2033 -734 -1999
rect -700 -2033 -694 -1999
rect -902 -2071 -694 -2033
rect -902 -2105 -896 -2071
rect -862 -2105 -815 -2071
rect -781 -2105 -734 -2071
rect -700 -2105 -694 -2071
rect -902 -2143 -694 -2105
rect -902 -2177 -896 -2143
rect -862 -2177 -815 -2143
rect -781 -2177 -734 -2143
rect -700 -2177 -694 -2143
rect -902 -2215 -694 -2177
rect -902 -2249 -896 -2215
rect -862 -2249 -815 -2215
rect -781 -2249 -734 -2215
rect -700 -2249 -694 -2215
rect -902 -2287 -694 -2249
rect -902 -2321 -896 -2287
rect -862 -2321 -815 -2287
rect -781 -2321 -734 -2287
rect -700 -2321 -694 -2287
rect -902 -2359 -694 -2321
rect -902 -2393 -896 -2359
rect -862 -2393 -815 -2359
rect -781 -2393 -734 -2359
rect -700 -2393 -694 -2359
rect -902 -2431 -694 -2393
rect -902 -2465 -896 -2431
rect -862 -2465 -815 -2431
rect -781 -2465 -734 -2431
rect -700 -2465 -694 -2431
rect -902 -2503 -694 -2465
rect -902 -2537 -896 -2503
rect -862 -2537 -815 -2503
rect -781 -2537 -734 -2503
rect -700 -2537 -694 -2503
rect -902 -2575 -694 -2537
rect -902 -2609 -896 -2575
rect -862 -2609 -815 -2575
rect -781 -2609 -734 -2575
rect -700 -2609 -694 -2575
rect -902 -2647 -694 -2609
rect -902 -2681 -896 -2647
rect -862 -2681 -815 -2647
rect -781 -2681 -734 -2647
rect -700 -2681 -694 -2647
rect -902 -2719 -694 -2681
rect -902 -2753 -896 -2719
rect -862 -2753 -815 -2719
rect -781 -2753 -734 -2719
rect -700 -2753 -694 -2719
rect -902 -2791 -694 -2753
rect -902 -2825 -896 -2791
rect -862 -2825 -815 -2791
rect -781 -2825 -734 -2791
rect -700 -2825 -694 -2791
rect -902 -2863 -694 -2825
rect -902 -2897 -896 -2863
rect -862 -2897 -815 -2863
rect -781 -2897 -734 -2863
rect -700 -2897 -694 -2863
rect -902 -2935 -694 -2897
rect -902 -2969 -896 -2935
rect -862 -2969 -815 -2935
rect -781 -2969 -734 -2935
rect -700 -2969 -694 -2935
rect -902 -3007 -694 -2969
rect -902 -3041 -896 -3007
rect -862 -3041 -815 -3007
rect -781 -3041 -734 -3007
rect -700 -3041 -694 -3007
rect -902 -3079 -694 -3041
rect -902 -3113 -896 -3079
rect -862 -3113 -815 -3079
rect -781 -3113 -734 -3079
rect -700 -3113 -694 -3079
rect -902 -3151 -694 -3113
rect -902 -3185 -896 -3151
rect -862 -3185 -815 -3151
rect -781 -3185 -734 -3151
rect -700 -3185 -694 -3151
rect -902 -3223 -694 -3185
rect -902 -3257 -896 -3223
rect -862 -3257 -815 -3223
rect -781 -3257 -734 -3223
rect -700 -3257 -694 -3223
rect -902 -3295 -694 -3257
rect -902 -3329 -896 -3295
rect -862 -3329 -815 -3295
rect -781 -3329 -734 -3295
rect -700 -3329 -694 -3295
rect -902 -3367 -694 -3329
rect -902 -3401 -896 -3367
rect -862 -3401 -815 -3367
rect -781 -3401 -734 -3367
rect -700 -3401 -694 -3367
rect -902 -3439 -694 -3401
rect -902 -3473 -896 -3439
rect -862 -3473 -815 -3439
rect -781 -3473 -734 -3439
rect -700 -3473 -694 -3439
rect -902 -3511 -694 -3473
rect -902 -3545 -896 -3511
rect -862 -3545 -815 -3511
rect -781 -3545 -734 -3511
rect -700 -3545 -694 -3511
rect -902 -3583 -694 -3545
rect -902 -3617 -896 -3583
rect -862 -3617 -815 -3583
rect -781 -3617 -734 -3583
rect -700 -3617 -694 -3583
rect -902 -3655 -694 -3617
rect -902 -3689 -896 -3655
rect -862 -3689 -815 -3655
rect -781 -3689 -734 -3655
rect -700 -3689 -694 -3655
rect -902 -3727 -694 -3689
rect -902 -3761 -896 -3727
rect -862 -3761 -815 -3727
rect -781 -3761 -734 -3727
rect -700 -3761 -694 -3727
rect -902 -3799 -694 -3761
rect -902 -3833 -896 -3799
rect -862 -3833 -815 -3799
rect -781 -3833 -734 -3799
rect -700 -3833 -694 -3799
rect -902 -3871 -694 -3833
rect -902 -3905 -896 -3871
rect -862 -3905 -815 -3871
rect -781 -3905 -734 -3871
rect -700 -3905 -694 -3871
rect -902 -3943 -694 -3905
rect -902 -3977 -896 -3943
rect -862 -3977 -815 -3943
rect -781 -3977 -734 -3943
rect -700 -3977 -694 -3943
rect -902 -4015 -694 -3977
rect -902 -4049 -896 -4015
rect -862 -4049 -815 -4015
rect -781 -4049 -734 -4015
rect -700 -4049 -694 -4015
rect -902 -4087 -694 -4049
rect -902 -4121 -896 -4087
rect -862 -4121 -815 -4087
rect -781 -4121 -734 -4087
rect -700 -4121 -694 -4087
rect -902 -4159 -694 -4121
rect -902 -4193 -896 -4159
rect -862 -4193 -815 -4159
rect -781 -4193 -734 -4159
rect -700 -4193 -694 -4159
rect -902 -4231 -694 -4193
rect -902 -4265 -896 -4231
rect -862 -4265 -815 -4231
rect -781 -4265 -734 -4231
rect -700 -4265 -694 -4231
rect -902 -4303 -694 -4265
rect -902 -4337 -896 -4303
rect -862 -4337 -815 -4303
rect -781 -4337 -734 -4303
rect -700 -4337 -694 -4303
rect -902 -4375 -694 -4337
rect -902 -4409 -896 -4375
rect -862 -4409 -815 -4375
rect -781 -4409 -734 -4375
rect -700 -4409 -694 -4375
rect -902 -4447 -694 -4409
rect -902 -4481 -896 -4447
rect -862 -4481 -815 -4447
rect -781 -4481 -734 -4447
rect -700 -4481 -694 -4447
rect -902 -4519 -694 -4481
rect -902 -4553 -896 -4519
rect -862 -4553 -815 -4519
rect -781 -4553 -734 -4519
rect -700 -4553 -694 -4519
rect -902 -4591 -694 -4553
rect -902 -4625 -896 -4591
rect -862 -4625 -815 -4591
rect -781 -4625 -734 -4591
rect -700 -4625 -694 -4591
rect -902 -4663 -694 -4625
rect -902 -4697 -896 -4663
rect -862 -4697 -815 -4663
rect -781 -4697 -734 -4663
rect -700 -4697 -694 -4663
rect -902 -4735 -694 -4697
rect -902 -4769 -896 -4735
rect -862 -4769 -815 -4735
rect -781 -4769 -734 -4735
rect -700 -4769 -694 -4735
rect -902 -4807 -694 -4769
rect -902 -4841 -896 -4807
rect -862 -4841 -815 -4807
rect -781 -4841 -734 -4807
rect -700 -4841 -694 -4807
rect -902 -4879 -694 -4841
rect -902 -4913 -896 -4879
rect -862 -4913 -815 -4879
rect -781 -4913 -734 -4879
rect -700 -4913 -694 -4879
rect -902 -4951 -694 -4913
rect -902 -4985 -896 -4951
rect -862 -4985 -815 -4951
rect -781 -4985 -734 -4951
rect -700 -4985 -694 -4951
tri -1226 -5062 -1186 -5022 sw
tri -942 -5062 -902 -5022 se
rect -902 -5062 -694 -4985
tri -626 5000 -606 5020 se
rect -606 5000 -458 5020
tri -458 5000 -438 5020 sw
rect -626 4985 -438 5000
rect -626 -4985 -585 4985
rect -479 -4985 -438 4985
rect -626 -5000 -438 -4985
tri -626 -5020 -606 -5000 ne
rect -606 -5020 -458 -5000
tri -458 -5020 -438 -5000 nw
rect -370 4985 -162 5062
tri -162 5022 -122 5062 nw
tri 122 5022 162 5062 ne
rect -370 4951 -364 4985
rect -330 4951 -283 4985
rect -249 4951 -202 4985
rect -168 4951 -162 4985
rect -370 4913 -162 4951
rect -370 4879 -364 4913
rect -330 4879 -283 4913
rect -249 4879 -202 4913
rect -168 4879 -162 4913
rect -370 4841 -162 4879
rect -370 4807 -364 4841
rect -330 4807 -283 4841
rect -249 4807 -202 4841
rect -168 4807 -162 4841
rect -370 4769 -162 4807
rect -370 4735 -364 4769
rect -330 4735 -283 4769
rect -249 4735 -202 4769
rect -168 4735 -162 4769
rect -370 4697 -162 4735
rect -370 4663 -364 4697
rect -330 4663 -283 4697
rect -249 4663 -202 4697
rect -168 4663 -162 4697
rect -370 4625 -162 4663
rect -370 4591 -364 4625
rect -330 4591 -283 4625
rect -249 4591 -202 4625
rect -168 4591 -162 4625
rect -370 4553 -162 4591
rect -370 4519 -364 4553
rect -330 4519 -283 4553
rect -249 4519 -202 4553
rect -168 4519 -162 4553
rect -370 4481 -162 4519
rect -370 4447 -364 4481
rect -330 4447 -283 4481
rect -249 4447 -202 4481
rect -168 4447 -162 4481
rect -370 4409 -162 4447
rect -370 4375 -364 4409
rect -330 4375 -283 4409
rect -249 4375 -202 4409
rect -168 4375 -162 4409
rect -370 4337 -162 4375
rect -370 4303 -364 4337
rect -330 4303 -283 4337
rect -249 4303 -202 4337
rect -168 4303 -162 4337
rect -370 4265 -162 4303
rect -370 4231 -364 4265
rect -330 4231 -283 4265
rect -249 4231 -202 4265
rect -168 4231 -162 4265
rect -370 4193 -162 4231
rect -370 4159 -364 4193
rect -330 4159 -283 4193
rect -249 4159 -202 4193
rect -168 4159 -162 4193
rect -370 4121 -162 4159
rect -370 4087 -364 4121
rect -330 4087 -283 4121
rect -249 4087 -202 4121
rect -168 4087 -162 4121
rect -370 4049 -162 4087
rect -370 4015 -364 4049
rect -330 4015 -283 4049
rect -249 4015 -202 4049
rect -168 4015 -162 4049
rect -370 3977 -162 4015
rect -370 3943 -364 3977
rect -330 3943 -283 3977
rect -249 3943 -202 3977
rect -168 3943 -162 3977
rect -370 3905 -162 3943
rect -370 3871 -364 3905
rect -330 3871 -283 3905
rect -249 3871 -202 3905
rect -168 3871 -162 3905
rect -370 3833 -162 3871
rect -370 3799 -364 3833
rect -330 3799 -283 3833
rect -249 3799 -202 3833
rect -168 3799 -162 3833
rect -370 3761 -162 3799
rect -370 3727 -364 3761
rect -330 3727 -283 3761
rect -249 3727 -202 3761
rect -168 3727 -162 3761
rect -370 3689 -162 3727
rect -370 3655 -364 3689
rect -330 3655 -283 3689
rect -249 3655 -202 3689
rect -168 3655 -162 3689
rect -370 3617 -162 3655
rect -370 3583 -364 3617
rect -330 3583 -283 3617
rect -249 3583 -202 3617
rect -168 3583 -162 3617
rect -370 3545 -162 3583
rect -370 3511 -364 3545
rect -330 3511 -283 3545
rect -249 3511 -202 3545
rect -168 3511 -162 3545
rect -370 3473 -162 3511
rect -370 3439 -364 3473
rect -330 3439 -283 3473
rect -249 3439 -202 3473
rect -168 3439 -162 3473
rect -370 3401 -162 3439
rect -370 3367 -364 3401
rect -330 3367 -283 3401
rect -249 3367 -202 3401
rect -168 3367 -162 3401
rect -370 3329 -162 3367
rect -370 3295 -364 3329
rect -330 3295 -283 3329
rect -249 3295 -202 3329
rect -168 3295 -162 3329
rect -370 3257 -162 3295
rect -370 3223 -364 3257
rect -330 3223 -283 3257
rect -249 3223 -202 3257
rect -168 3223 -162 3257
rect -370 3185 -162 3223
rect -370 3151 -364 3185
rect -330 3151 -283 3185
rect -249 3151 -202 3185
rect -168 3151 -162 3185
rect -370 3113 -162 3151
rect -370 3079 -364 3113
rect -330 3079 -283 3113
rect -249 3079 -202 3113
rect -168 3079 -162 3113
rect -370 3041 -162 3079
rect -370 3007 -364 3041
rect -330 3007 -283 3041
rect -249 3007 -202 3041
rect -168 3007 -162 3041
rect -370 2969 -162 3007
rect -370 2935 -364 2969
rect -330 2935 -283 2969
rect -249 2935 -202 2969
rect -168 2935 -162 2969
rect -370 2897 -162 2935
rect -370 2863 -364 2897
rect -330 2863 -283 2897
rect -249 2863 -202 2897
rect -168 2863 -162 2897
rect -370 2825 -162 2863
rect -370 2791 -364 2825
rect -330 2791 -283 2825
rect -249 2791 -202 2825
rect -168 2791 -162 2825
rect -370 2753 -162 2791
rect -370 2719 -364 2753
rect -330 2719 -283 2753
rect -249 2719 -202 2753
rect -168 2719 -162 2753
rect -370 2681 -162 2719
rect -370 2647 -364 2681
rect -330 2647 -283 2681
rect -249 2647 -202 2681
rect -168 2647 -162 2681
rect -370 2609 -162 2647
rect -370 2575 -364 2609
rect -330 2575 -283 2609
rect -249 2575 -202 2609
rect -168 2575 -162 2609
rect -370 2537 -162 2575
rect -370 2503 -364 2537
rect -330 2503 -283 2537
rect -249 2503 -202 2537
rect -168 2503 -162 2537
rect -370 2465 -162 2503
rect -370 2431 -364 2465
rect -330 2431 -283 2465
rect -249 2431 -202 2465
rect -168 2431 -162 2465
rect -370 2393 -162 2431
rect -370 2359 -364 2393
rect -330 2359 -283 2393
rect -249 2359 -202 2393
rect -168 2359 -162 2393
rect -370 2321 -162 2359
rect -370 2287 -364 2321
rect -330 2287 -283 2321
rect -249 2287 -202 2321
rect -168 2287 -162 2321
rect -370 2249 -162 2287
rect -370 2215 -364 2249
rect -330 2215 -283 2249
rect -249 2215 -202 2249
rect -168 2215 -162 2249
rect -370 2177 -162 2215
rect -370 2143 -364 2177
rect -330 2143 -283 2177
rect -249 2143 -202 2177
rect -168 2143 -162 2177
rect -370 2105 -162 2143
rect -370 2071 -364 2105
rect -330 2071 -283 2105
rect -249 2071 -202 2105
rect -168 2071 -162 2105
rect -370 2033 -162 2071
rect -370 1999 -364 2033
rect -330 1999 -283 2033
rect -249 1999 -202 2033
rect -168 1999 -162 2033
rect -370 1961 -162 1999
rect -370 1927 -364 1961
rect -330 1927 -283 1961
rect -249 1927 -202 1961
rect -168 1927 -162 1961
rect -370 1889 -162 1927
rect -370 1855 -364 1889
rect -330 1855 -283 1889
rect -249 1855 -202 1889
rect -168 1855 -162 1889
rect -370 1817 -162 1855
rect -370 1783 -364 1817
rect -330 1783 -283 1817
rect -249 1783 -202 1817
rect -168 1783 -162 1817
rect -370 1745 -162 1783
rect -370 1711 -364 1745
rect -330 1711 -283 1745
rect -249 1711 -202 1745
rect -168 1711 -162 1745
rect -370 1673 -162 1711
rect -370 1639 -364 1673
rect -330 1639 -283 1673
rect -249 1639 -202 1673
rect -168 1639 -162 1673
rect -370 1601 -162 1639
rect -370 1567 -364 1601
rect -330 1567 -283 1601
rect -249 1567 -202 1601
rect -168 1567 -162 1601
rect -370 1529 -162 1567
rect -370 1495 -364 1529
rect -330 1495 -283 1529
rect -249 1495 -202 1529
rect -168 1495 -162 1529
rect -370 1457 -162 1495
rect -370 1423 -364 1457
rect -330 1423 -283 1457
rect -249 1423 -202 1457
rect -168 1423 -162 1457
rect -370 1385 -162 1423
rect -370 1351 -364 1385
rect -330 1351 -283 1385
rect -249 1351 -202 1385
rect -168 1351 -162 1385
rect -370 1313 -162 1351
rect -370 1279 -364 1313
rect -330 1279 -283 1313
rect -249 1279 -202 1313
rect -168 1279 -162 1313
rect -370 1241 -162 1279
rect -370 1207 -364 1241
rect -330 1207 -283 1241
rect -249 1207 -202 1241
rect -168 1207 -162 1241
rect -370 1169 -162 1207
rect -370 1135 -364 1169
rect -330 1135 -283 1169
rect -249 1135 -202 1169
rect -168 1135 -162 1169
rect -370 1097 -162 1135
rect -370 1063 -364 1097
rect -330 1063 -283 1097
rect -249 1063 -202 1097
rect -168 1063 -162 1097
rect -370 1025 -162 1063
rect -370 991 -364 1025
rect -330 991 -283 1025
rect -249 991 -202 1025
rect -168 991 -162 1025
rect -370 953 -162 991
rect -370 919 -364 953
rect -330 919 -283 953
rect -249 919 -202 953
rect -168 919 -162 953
rect -370 881 -162 919
rect -370 847 -364 881
rect -330 847 -283 881
rect -249 847 -202 881
rect -168 847 -162 881
rect -370 809 -162 847
rect -370 775 -364 809
rect -330 775 -283 809
rect -249 775 -202 809
rect -168 775 -162 809
rect -370 737 -162 775
rect -370 703 -364 737
rect -330 703 -283 737
rect -249 703 -202 737
rect -168 703 -162 737
rect -370 665 -162 703
rect -370 631 -364 665
rect -330 631 -283 665
rect -249 631 -202 665
rect -168 631 -162 665
rect -370 593 -162 631
rect -370 559 -364 593
rect -330 559 -283 593
rect -249 559 -202 593
rect -168 559 -162 593
rect -370 521 -162 559
rect -370 487 -364 521
rect -330 487 -283 521
rect -249 487 -202 521
rect -168 487 -162 521
rect -370 449 -162 487
rect -370 415 -364 449
rect -330 415 -283 449
rect -249 415 -202 449
rect -168 415 -162 449
rect -370 377 -162 415
rect -370 343 -364 377
rect -330 343 -283 377
rect -249 343 -202 377
rect -168 343 -162 377
rect -370 305 -162 343
rect -370 271 -364 305
rect -330 271 -283 305
rect -249 271 -202 305
rect -168 271 -162 305
rect -370 233 -162 271
rect -370 199 -364 233
rect -330 199 -283 233
rect -249 199 -202 233
rect -168 199 -162 233
rect -370 161 -162 199
rect -370 127 -364 161
rect -330 127 -283 161
rect -249 127 -202 161
rect -168 127 -162 161
rect -370 89 -162 127
rect -370 55 -364 89
rect -330 55 -283 89
rect -249 55 -202 89
rect -168 55 -162 89
rect -370 17 -162 55
rect -370 -17 -364 17
rect -330 -17 -283 17
rect -249 -17 -202 17
rect -168 -17 -162 17
rect -370 -55 -162 -17
rect -370 -89 -364 -55
rect -330 -89 -283 -55
rect -249 -89 -202 -55
rect -168 -89 -162 -55
rect -370 -127 -162 -89
rect -370 -161 -364 -127
rect -330 -161 -283 -127
rect -249 -161 -202 -127
rect -168 -161 -162 -127
rect -370 -199 -162 -161
rect -370 -233 -364 -199
rect -330 -233 -283 -199
rect -249 -233 -202 -199
rect -168 -233 -162 -199
rect -370 -271 -162 -233
rect -370 -305 -364 -271
rect -330 -305 -283 -271
rect -249 -305 -202 -271
rect -168 -305 -162 -271
rect -370 -343 -162 -305
rect -370 -377 -364 -343
rect -330 -377 -283 -343
rect -249 -377 -202 -343
rect -168 -377 -162 -343
rect -370 -415 -162 -377
rect -370 -449 -364 -415
rect -330 -449 -283 -415
rect -249 -449 -202 -415
rect -168 -449 -162 -415
rect -370 -487 -162 -449
rect -370 -521 -364 -487
rect -330 -521 -283 -487
rect -249 -521 -202 -487
rect -168 -521 -162 -487
rect -370 -559 -162 -521
rect -370 -593 -364 -559
rect -330 -593 -283 -559
rect -249 -593 -202 -559
rect -168 -593 -162 -559
rect -370 -631 -162 -593
rect -370 -665 -364 -631
rect -330 -665 -283 -631
rect -249 -665 -202 -631
rect -168 -665 -162 -631
rect -370 -703 -162 -665
rect -370 -737 -364 -703
rect -330 -737 -283 -703
rect -249 -737 -202 -703
rect -168 -737 -162 -703
rect -370 -775 -162 -737
rect -370 -809 -364 -775
rect -330 -809 -283 -775
rect -249 -809 -202 -775
rect -168 -809 -162 -775
rect -370 -847 -162 -809
rect -370 -881 -364 -847
rect -330 -881 -283 -847
rect -249 -881 -202 -847
rect -168 -881 -162 -847
rect -370 -919 -162 -881
rect -370 -953 -364 -919
rect -330 -953 -283 -919
rect -249 -953 -202 -919
rect -168 -953 -162 -919
rect -370 -991 -162 -953
rect -370 -1025 -364 -991
rect -330 -1025 -283 -991
rect -249 -1025 -202 -991
rect -168 -1025 -162 -991
rect -370 -1063 -162 -1025
rect -370 -1097 -364 -1063
rect -330 -1097 -283 -1063
rect -249 -1097 -202 -1063
rect -168 -1097 -162 -1063
rect -370 -1135 -162 -1097
rect -370 -1169 -364 -1135
rect -330 -1169 -283 -1135
rect -249 -1169 -202 -1135
rect -168 -1169 -162 -1135
rect -370 -1207 -162 -1169
rect -370 -1241 -364 -1207
rect -330 -1241 -283 -1207
rect -249 -1241 -202 -1207
rect -168 -1241 -162 -1207
rect -370 -1279 -162 -1241
rect -370 -1313 -364 -1279
rect -330 -1313 -283 -1279
rect -249 -1313 -202 -1279
rect -168 -1313 -162 -1279
rect -370 -1351 -162 -1313
rect -370 -1385 -364 -1351
rect -330 -1385 -283 -1351
rect -249 -1385 -202 -1351
rect -168 -1385 -162 -1351
rect -370 -1423 -162 -1385
rect -370 -1457 -364 -1423
rect -330 -1457 -283 -1423
rect -249 -1457 -202 -1423
rect -168 -1457 -162 -1423
rect -370 -1495 -162 -1457
rect -370 -1529 -364 -1495
rect -330 -1529 -283 -1495
rect -249 -1529 -202 -1495
rect -168 -1529 -162 -1495
rect -370 -1567 -162 -1529
rect -370 -1601 -364 -1567
rect -330 -1601 -283 -1567
rect -249 -1601 -202 -1567
rect -168 -1601 -162 -1567
rect -370 -1639 -162 -1601
rect -370 -1673 -364 -1639
rect -330 -1673 -283 -1639
rect -249 -1673 -202 -1639
rect -168 -1673 -162 -1639
rect -370 -1711 -162 -1673
rect -370 -1745 -364 -1711
rect -330 -1745 -283 -1711
rect -249 -1745 -202 -1711
rect -168 -1745 -162 -1711
rect -370 -1783 -162 -1745
rect -370 -1817 -364 -1783
rect -330 -1817 -283 -1783
rect -249 -1817 -202 -1783
rect -168 -1817 -162 -1783
rect -370 -1855 -162 -1817
rect -370 -1889 -364 -1855
rect -330 -1889 -283 -1855
rect -249 -1889 -202 -1855
rect -168 -1889 -162 -1855
rect -370 -1927 -162 -1889
rect -370 -1961 -364 -1927
rect -330 -1961 -283 -1927
rect -249 -1961 -202 -1927
rect -168 -1961 -162 -1927
rect -370 -1999 -162 -1961
rect -370 -2033 -364 -1999
rect -330 -2033 -283 -1999
rect -249 -2033 -202 -1999
rect -168 -2033 -162 -1999
rect -370 -2071 -162 -2033
rect -370 -2105 -364 -2071
rect -330 -2105 -283 -2071
rect -249 -2105 -202 -2071
rect -168 -2105 -162 -2071
rect -370 -2143 -162 -2105
rect -370 -2177 -364 -2143
rect -330 -2177 -283 -2143
rect -249 -2177 -202 -2143
rect -168 -2177 -162 -2143
rect -370 -2215 -162 -2177
rect -370 -2249 -364 -2215
rect -330 -2249 -283 -2215
rect -249 -2249 -202 -2215
rect -168 -2249 -162 -2215
rect -370 -2287 -162 -2249
rect -370 -2321 -364 -2287
rect -330 -2321 -283 -2287
rect -249 -2321 -202 -2287
rect -168 -2321 -162 -2287
rect -370 -2359 -162 -2321
rect -370 -2393 -364 -2359
rect -330 -2393 -283 -2359
rect -249 -2393 -202 -2359
rect -168 -2393 -162 -2359
rect -370 -2431 -162 -2393
rect -370 -2465 -364 -2431
rect -330 -2465 -283 -2431
rect -249 -2465 -202 -2431
rect -168 -2465 -162 -2431
rect -370 -2503 -162 -2465
rect -370 -2537 -364 -2503
rect -330 -2537 -283 -2503
rect -249 -2537 -202 -2503
rect -168 -2537 -162 -2503
rect -370 -2575 -162 -2537
rect -370 -2609 -364 -2575
rect -330 -2609 -283 -2575
rect -249 -2609 -202 -2575
rect -168 -2609 -162 -2575
rect -370 -2647 -162 -2609
rect -370 -2681 -364 -2647
rect -330 -2681 -283 -2647
rect -249 -2681 -202 -2647
rect -168 -2681 -162 -2647
rect -370 -2719 -162 -2681
rect -370 -2753 -364 -2719
rect -330 -2753 -283 -2719
rect -249 -2753 -202 -2719
rect -168 -2753 -162 -2719
rect -370 -2791 -162 -2753
rect -370 -2825 -364 -2791
rect -330 -2825 -283 -2791
rect -249 -2825 -202 -2791
rect -168 -2825 -162 -2791
rect -370 -2863 -162 -2825
rect -370 -2897 -364 -2863
rect -330 -2897 -283 -2863
rect -249 -2897 -202 -2863
rect -168 -2897 -162 -2863
rect -370 -2935 -162 -2897
rect -370 -2969 -364 -2935
rect -330 -2969 -283 -2935
rect -249 -2969 -202 -2935
rect -168 -2969 -162 -2935
rect -370 -3007 -162 -2969
rect -370 -3041 -364 -3007
rect -330 -3041 -283 -3007
rect -249 -3041 -202 -3007
rect -168 -3041 -162 -3007
rect -370 -3079 -162 -3041
rect -370 -3113 -364 -3079
rect -330 -3113 -283 -3079
rect -249 -3113 -202 -3079
rect -168 -3113 -162 -3079
rect -370 -3151 -162 -3113
rect -370 -3185 -364 -3151
rect -330 -3185 -283 -3151
rect -249 -3185 -202 -3151
rect -168 -3185 -162 -3151
rect -370 -3223 -162 -3185
rect -370 -3257 -364 -3223
rect -330 -3257 -283 -3223
rect -249 -3257 -202 -3223
rect -168 -3257 -162 -3223
rect -370 -3295 -162 -3257
rect -370 -3329 -364 -3295
rect -330 -3329 -283 -3295
rect -249 -3329 -202 -3295
rect -168 -3329 -162 -3295
rect -370 -3367 -162 -3329
rect -370 -3401 -364 -3367
rect -330 -3401 -283 -3367
rect -249 -3401 -202 -3367
rect -168 -3401 -162 -3367
rect -370 -3439 -162 -3401
rect -370 -3473 -364 -3439
rect -330 -3473 -283 -3439
rect -249 -3473 -202 -3439
rect -168 -3473 -162 -3439
rect -370 -3511 -162 -3473
rect -370 -3545 -364 -3511
rect -330 -3545 -283 -3511
rect -249 -3545 -202 -3511
rect -168 -3545 -162 -3511
rect -370 -3583 -162 -3545
rect -370 -3617 -364 -3583
rect -330 -3617 -283 -3583
rect -249 -3617 -202 -3583
rect -168 -3617 -162 -3583
rect -370 -3655 -162 -3617
rect -370 -3689 -364 -3655
rect -330 -3689 -283 -3655
rect -249 -3689 -202 -3655
rect -168 -3689 -162 -3655
rect -370 -3727 -162 -3689
rect -370 -3761 -364 -3727
rect -330 -3761 -283 -3727
rect -249 -3761 -202 -3727
rect -168 -3761 -162 -3727
rect -370 -3799 -162 -3761
rect -370 -3833 -364 -3799
rect -330 -3833 -283 -3799
rect -249 -3833 -202 -3799
rect -168 -3833 -162 -3799
rect -370 -3871 -162 -3833
rect -370 -3905 -364 -3871
rect -330 -3905 -283 -3871
rect -249 -3905 -202 -3871
rect -168 -3905 -162 -3871
rect -370 -3943 -162 -3905
rect -370 -3977 -364 -3943
rect -330 -3977 -283 -3943
rect -249 -3977 -202 -3943
rect -168 -3977 -162 -3943
rect -370 -4015 -162 -3977
rect -370 -4049 -364 -4015
rect -330 -4049 -283 -4015
rect -249 -4049 -202 -4015
rect -168 -4049 -162 -4015
rect -370 -4087 -162 -4049
rect -370 -4121 -364 -4087
rect -330 -4121 -283 -4087
rect -249 -4121 -202 -4087
rect -168 -4121 -162 -4087
rect -370 -4159 -162 -4121
rect -370 -4193 -364 -4159
rect -330 -4193 -283 -4159
rect -249 -4193 -202 -4159
rect -168 -4193 -162 -4159
rect -370 -4231 -162 -4193
rect -370 -4265 -364 -4231
rect -330 -4265 -283 -4231
rect -249 -4265 -202 -4231
rect -168 -4265 -162 -4231
rect -370 -4303 -162 -4265
rect -370 -4337 -364 -4303
rect -330 -4337 -283 -4303
rect -249 -4337 -202 -4303
rect -168 -4337 -162 -4303
rect -370 -4375 -162 -4337
rect -370 -4409 -364 -4375
rect -330 -4409 -283 -4375
rect -249 -4409 -202 -4375
rect -168 -4409 -162 -4375
rect -370 -4447 -162 -4409
rect -370 -4481 -364 -4447
rect -330 -4481 -283 -4447
rect -249 -4481 -202 -4447
rect -168 -4481 -162 -4447
rect -370 -4519 -162 -4481
rect -370 -4553 -364 -4519
rect -330 -4553 -283 -4519
rect -249 -4553 -202 -4519
rect -168 -4553 -162 -4519
rect -370 -4591 -162 -4553
rect -370 -4625 -364 -4591
rect -330 -4625 -283 -4591
rect -249 -4625 -202 -4591
rect -168 -4625 -162 -4591
rect -370 -4663 -162 -4625
rect -370 -4697 -364 -4663
rect -330 -4697 -283 -4663
rect -249 -4697 -202 -4663
rect -168 -4697 -162 -4663
rect -370 -4735 -162 -4697
rect -370 -4769 -364 -4735
rect -330 -4769 -283 -4735
rect -249 -4769 -202 -4735
rect -168 -4769 -162 -4735
rect -370 -4807 -162 -4769
rect -370 -4841 -364 -4807
rect -330 -4841 -283 -4807
rect -249 -4841 -202 -4807
rect -168 -4841 -162 -4807
rect -370 -4879 -162 -4841
rect -370 -4913 -364 -4879
rect -330 -4913 -283 -4879
rect -249 -4913 -202 -4879
rect -168 -4913 -162 -4879
rect -370 -4951 -162 -4913
rect -370 -4985 -364 -4951
rect -330 -4985 -283 -4951
rect -249 -4985 -202 -4951
rect -168 -4985 -162 -4951
tri -694 -5062 -654 -5022 sw
tri -410 -5062 -370 -5022 se
rect -370 -5062 -162 -4985
tri -94 5000 -74 5020 se
rect -74 5000 74 5020
tri 74 5000 94 5020 sw
rect -94 4985 94 5000
rect -94 -4985 -53 4985
rect 53 -4985 94 4985
rect -94 -5000 94 -4985
tri -94 -5020 -74 -5000 ne
rect -74 -5020 74 -5000
tri 74 -5020 94 -5000 nw
rect 162 4985 370 5062
tri 370 5022 410 5062 nw
tri 654 5022 694 5062 ne
rect 162 4951 168 4985
rect 202 4951 249 4985
rect 283 4951 330 4985
rect 364 4951 370 4985
rect 162 4913 370 4951
rect 162 4879 168 4913
rect 202 4879 249 4913
rect 283 4879 330 4913
rect 364 4879 370 4913
rect 162 4841 370 4879
rect 162 4807 168 4841
rect 202 4807 249 4841
rect 283 4807 330 4841
rect 364 4807 370 4841
rect 162 4769 370 4807
rect 162 4735 168 4769
rect 202 4735 249 4769
rect 283 4735 330 4769
rect 364 4735 370 4769
rect 162 4697 370 4735
rect 162 4663 168 4697
rect 202 4663 249 4697
rect 283 4663 330 4697
rect 364 4663 370 4697
rect 162 4625 370 4663
rect 162 4591 168 4625
rect 202 4591 249 4625
rect 283 4591 330 4625
rect 364 4591 370 4625
rect 162 4553 370 4591
rect 162 4519 168 4553
rect 202 4519 249 4553
rect 283 4519 330 4553
rect 364 4519 370 4553
rect 162 4481 370 4519
rect 162 4447 168 4481
rect 202 4447 249 4481
rect 283 4447 330 4481
rect 364 4447 370 4481
rect 162 4409 370 4447
rect 162 4375 168 4409
rect 202 4375 249 4409
rect 283 4375 330 4409
rect 364 4375 370 4409
rect 162 4337 370 4375
rect 162 4303 168 4337
rect 202 4303 249 4337
rect 283 4303 330 4337
rect 364 4303 370 4337
rect 162 4265 370 4303
rect 162 4231 168 4265
rect 202 4231 249 4265
rect 283 4231 330 4265
rect 364 4231 370 4265
rect 162 4193 370 4231
rect 162 4159 168 4193
rect 202 4159 249 4193
rect 283 4159 330 4193
rect 364 4159 370 4193
rect 162 4121 370 4159
rect 162 4087 168 4121
rect 202 4087 249 4121
rect 283 4087 330 4121
rect 364 4087 370 4121
rect 162 4049 370 4087
rect 162 4015 168 4049
rect 202 4015 249 4049
rect 283 4015 330 4049
rect 364 4015 370 4049
rect 162 3977 370 4015
rect 162 3943 168 3977
rect 202 3943 249 3977
rect 283 3943 330 3977
rect 364 3943 370 3977
rect 162 3905 370 3943
rect 162 3871 168 3905
rect 202 3871 249 3905
rect 283 3871 330 3905
rect 364 3871 370 3905
rect 162 3833 370 3871
rect 162 3799 168 3833
rect 202 3799 249 3833
rect 283 3799 330 3833
rect 364 3799 370 3833
rect 162 3761 370 3799
rect 162 3727 168 3761
rect 202 3727 249 3761
rect 283 3727 330 3761
rect 364 3727 370 3761
rect 162 3689 370 3727
rect 162 3655 168 3689
rect 202 3655 249 3689
rect 283 3655 330 3689
rect 364 3655 370 3689
rect 162 3617 370 3655
rect 162 3583 168 3617
rect 202 3583 249 3617
rect 283 3583 330 3617
rect 364 3583 370 3617
rect 162 3545 370 3583
rect 162 3511 168 3545
rect 202 3511 249 3545
rect 283 3511 330 3545
rect 364 3511 370 3545
rect 162 3473 370 3511
rect 162 3439 168 3473
rect 202 3439 249 3473
rect 283 3439 330 3473
rect 364 3439 370 3473
rect 162 3401 370 3439
rect 162 3367 168 3401
rect 202 3367 249 3401
rect 283 3367 330 3401
rect 364 3367 370 3401
rect 162 3329 370 3367
rect 162 3295 168 3329
rect 202 3295 249 3329
rect 283 3295 330 3329
rect 364 3295 370 3329
rect 162 3257 370 3295
rect 162 3223 168 3257
rect 202 3223 249 3257
rect 283 3223 330 3257
rect 364 3223 370 3257
rect 162 3185 370 3223
rect 162 3151 168 3185
rect 202 3151 249 3185
rect 283 3151 330 3185
rect 364 3151 370 3185
rect 162 3113 370 3151
rect 162 3079 168 3113
rect 202 3079 249 3113
rect 283 3079 330 3113
rect 364 3079 370 3113
rect 162 3041 370 3079
rect 162 3007 168 3041
rect 202 3007 249 3041
rect 283 3007 330 3041
rect 364 3007 370 3041
rect 162 2969 370 3007
rect 162 2935 168 2969
rect 202 2935 249 2969
rect 283 2935 330 2969
rect 364 2935 370 2969
rect 162 2897 370 2935
rect 162 2863 168 2897
rect 202 2863 249 2897
rect 283 2863 330 2897
rect 364 2863 370 2897
rect 162 2825 370 2863
rect 162 2791 168 2825
rect 202 2791 249 2825
rect 283 2791 330 2825
rect 364 2791 370 2825
rect 162 2753 370 2791
rect 162 2719 168 2753
rect 202 2719 249 2753
rect 283 2719 330 2753
rect 364 2719 370 2753
rect 162 2681 370 2719
rect 162 2647 168 2681
rect 202 2647 249 2681
rect 283 2647 330 2681
rect 364 2647 370 2681
rect 162 2609 370 2647
rect 162 2575 168 2609
rect 202 2575 249 2609
rect 283 2575 330 2609
rect 364 2575 370 2609
rect 162 2537 370 2575
rect 162 2503 168 2537
rect 202 2503 249 2537
rect 283 2503 330 2537
rect 364 2503 370 2537
rect 162 2465 370 2503
rect 162 2431 168 2465
rect 202 2431 249 2465
rect 283 2431 330 2465
rect 364 2431 370 2465
rect 162 2393 370 2431
rect 162 2359 168 2393
rect 202 2359 249 2393
rect 283 2359 330 2393
rect 364 2359 370 2393
rect 162 2321 370 2359
rect 162 2287 168 2321
rect 202 2287 249 2321
rect 283 2287 330 2321
rect 364 2287 370 2321
rect 162 2249 370 2287
rect 162 2215 168 2249
rect 202 2215 249 2249
rect 283 2215 330 2249
rect 364 2215 370 2249
rect 162 2177 370 2215
rect 162 2143 168 2177
rect 202 2143 249 2177
rect 283 2143 330 2177
rect 364 2143 370 2177
rect 162 2105 370 2143
rect 162 2071 168 2105
rect 202 2071 249 2105
rect 283 2071 330 2105
rect 364 2071 370 2105
rect 162 2033 370 2071
rect 162 1999 168 2033
rect 202 1999 249 2033
rect 283 1999 330 2033
rect 364 1999 370 2033
rect 162 1961 370 1999
rect 162 1927 168 1961
rect 202 1927 249 1961
rect 283 1927 330 1961
rect 364 1927 370 1961
rect 162 1889 370 1927
rect 162 1855 168 1889
rect 202 1855 249 1889
rect 283 1855 330 1889
rect 364 1855 370 1889
rect 162 1817 370 1855
rect 162 1783 168 1817
rect 202 1783 249 1817
rect 283 1783 330 1817
rect 364 1783 370 1817
rect 162 1745 370 1783
rect 162 1711 168 1745
rect 202 1711 249 1745
rect 283 1711 330 1745
rect 364 1711 370 1745
rect 162 1673 370 1711
rect 162 1639 168 1673
rect 202 1639 249 1673
rect 283 1639 330 1673
rect 364 1639 370 1673
rect 162 1601 370 1639
rect 162 1567 168 1601
rect 202 1567 249 1601
rect 283 1567 330 1601
rect 364 1567 370 1601
rect 162 1529 370 1567
rect 162 1495 168 1529
rect 202 1495 249 1529
rect 283 1495 330 1529
rect 364 1495 370 1529
rect 162 1457 370 1495
rect 162 1423 168 1457
rect 202 1423 249 1457
rect 283 1423 330 1457
rect 364 1423 370 1457
rect 162 1385 370 1423
rect 162 1351 168 1385
rect 202 1351 249 1385
rect 283 1351 330 1385
rect 364 1351 370 1385
rect 162 1313 370 1351
rect 162 1279 168 1313
rect 202 1279 249 1313
rect 283 1279 330 1313
rect 364 1279 370 1313
rect 162 1241 370 1279
rect 162 1207 168 1241
rect 202 1207 249 1241
rect 283 1207 330 1241
rect 364 1207 370 1241
rect 162 1169 370 1207
rect 162 1135 168 1169
rect 202 1135 249 1169
rect 283 1135 330 1169
rect 364 1135 370 1169
rect 162 1097 370 1135
rect 162 1063 168 1097
rect 202 1063 249 1097
rect 283 1063 330 1097
rect 364 1063 370 1097
rect 162 1025 370 1063
rect 162 991 168 1025
rect 202 991 249 1025
rect 283 991 330 1025
rect 364 991 370 1025
rect 162 953 370 991
rect 162 919 168 953
rect 202 919 249 953
rect 283 919 330 953
rect 364 919 370 953
rect 162 881 370 919
rect 162 847 168 881
rect 202 847 249 881
rect 283 847 330 881
rect 364 847 370 881
rect 162 809 370 847
rect 162 775 168 809
rect 202 775 249 809
rect 283 775 330 809
rect 364 775 370 809
rect 162 737 370 775
rect 162 703 168 737
rect 202 703 249 737
rect 283 703 330 737
rect 364 703 370 737
rect 162 665 370 703
rect 162 631 168 665
rect 202 631 249 665
rect 283 631 330 665
rect 364 631 370 665
rect 162 593 370 631
rect 162 559 168 593
rect 202 559 249 593
rect 283 559 330 593
rect 364 559 370 593
rect 162 521 370 559
rect 162 487 168 521
rect 202 487 249 521
rect 283 487 330 521
rect 364 487 370 521
rect 162 449 370 487
rect 162 415 168 449
rect 202 415 249 449
rect 283 415 330 449
rect 364 415 370 449
rect 162 377 370 415
rect 162 343 168 377
rect 202 343 249 377
rect 283 343 330 377
rect 364 343 370 377
rect 162 305 370 343
rect 162 271 168 305
rect 202 271 249 305
rect 283 271 330 305
rect 364 271 370 305
rect 162 233 370 271
rect 162 199 168 233
rect 202 199 249 233
rect 283 199 330 233
rect 364 199 370 233
rect 162 161 370 199
rect 162 127 168 161
rect 202 127 249 161
rect 283 127 330 161
rect 364 127 370 161
rect 162 89 370 127
rect 162 55 168 89
rect 202 55 249 89
rect 283 55 330 89
rect 364 55 370 89
rect 162 17 370 55
rect 162 -17 168 17
rect 202 -17 249 17
rect 283 -17 330 17
rect 364 -17 370 17
rect 162 -55 370 -17
rect 162 -89 168 -55
rect 202 -89 249 -55
rect 283 -89 330 -55
rect 364 -89 370 -55
rect 162 -127 370 -89
rect 162 -161 168 -127
rect 202 -161 249 -127
rect 283 -161 330 -127
rect 364 -161 370 -127
rect 162 -199 370 -161
rect 162 -233 168 -199
rect 202 -233 249 -199
rect 283 -233 330 -199
rect 364 -233 370 -199
rect 162 -271 370 -233
rect 162 -305 168 -271
rect 202 -305 249 -271
rect 283 -305 330 -271
rect 364 -305 370 -271
rect 162 -343 370 -305
rect 162 -377 168 -343
rect 202 -377 249 -343
rect 283 -377 330 -343
rect 364 -377 370 -343
rect 162 -415 370 -377
rect 162 -449 168 -415
rect 202 -449 249 -415
rect 283 -449 330 -415
rect 364 -449 370 -415
rect 162 -487 370 -449
rect 162 -521 168 -487
rect 202 -521 249 -487
rect 283 -521 330 -487
rect 364 -521 370 -487
rect 162 -559 370 -521
rect 162 -593 168 -559
rect 202 -593 249 -559
rect 283 -593 330 -559
rect 364 -593 370 -559
rect 162 -631 370 -593
rect 162 -665 168 -631
rect 202 -665 249 -631
rect 283 -665 330 -631
rect 364 -665 370 -631
rect 162 -703 370 -665
rect 162 -737 168 -703
rect 202 -737 249 -703
rect 283 -737 330 -703
rect 364 -737 370 -703
rect 162 -775 370 -737
rect 162 -809 168 -775
rect 202 -809 249 -775
rect 283 -809 330 -775
rect 364 -809 370 -775
rect 162 -847 370 -809
rect 162 -881 168 -847
rect 202 -881 249 -847
rect 283 -881 330 -847
rect 364 -881 370 -847
rect 162 -919 370 -881
rect 162 -953 168 -919
rect 202 -953 249 -919
rect 283 -953 330 -919
rect 364 -953 370 -919
rect 162 -991 370 -953
rect 162 -1025 168 -991
rect 202 -1025 249 -991
rect 283 -1025 330 -991
rect 364 -1025 370 -991
rect 162 -1063 370 -1025
rect 162 -1097 168 -1063
rect 202 -1097 249 -1063
rect 283 -1097 330 -1063
rect 364 -1097 370 -1063
rect 162 -1135 370 -1097
rect 162 -1169 168 -1135
rect 202 -1169 249 -1135
rect 283 -1169 330 -1135
rect 364 -1169 370 -1135
rect 162 -1207 370 -1169
rect 162 -1241 168 -1207
rect 202 -1241 249 -1207
rect 283 -1241 330 -1207
rect 364 -1241 370 -1207
rect 162 -1279 370 -1241
rect 162 -1313 168 -1279
rect 202 -1313 249 -1279
rect 283 -1313 330 -1279
rect 364 -1313 370 -1279
rect 162 -1351 370 -1313
rect 162 -1385 168 -1351
rect 202 -1385 249 -1351
rect 283 -1385 330 -1351
rect 364 -1385 370 -1351
rect 162 -1423 370 -1385
rect 162 -1457 168 -1423
rect 202 -1457 249 -1423
rect 283 -1457 330 -1423
rect 364 -1457 370 -1423
rect 162 -1495 370 -1457
rect 162 -1529 168 -1495
rect 202 -1529 249 -1495
rect 283 -1529 330 -1495
rect 364 -1529 370 -1495
rect 162 -1567 370 -1529
rect 162 -1601 168 -1567
rect 202 -1601 249 -1567
rect 283 -1601 330 -1567
rect 364 -1601 370 -1567
rect 162 -1639 370 -1601
rect 162 -1673 168 -1639
rect 202 -1673 249 -1639
rect 283 -1673 330 -1639
rect 364 -1673 370 -1639
rect 162 -1711 370 -1673
rect 162 -1745 168 -1711
rect 202 -1745 249 -1711
rect 283 -1745 330 -1711
rect 364 -1745 370 -1711
rect 162 -1783 370 -1745
rect 162 -1817 168 -1783
rect 202 -1817 249 -1783
rect 283 -1817 330 -1783
rect 364 -1817 370 -1783
rect 162 -1855 370 -1817
rect 162 -1889 168 -1855
rect 202 -1889 249 -1855
rect 283 -1889 330 -1855
rect 364 -1889 370 -1855
rect 162 -1927 370 -1889
rect 162 -1961 168 -1927
rect 202 -1961 249 -1927
rect 283 -1961 330 -1927
rect 364 -1961 370 -1927
rect 162 -1999 370 -1961
rect 162 -2033 168 -1999
rect 202 -2033 249 -1999
rect 283 -2033 330 -1999
rect 364 -2033 370 -1999
rect 162 -2071 370 -2033
rect 162 -2105 168 -2071
rect 202 -2105 249 -2071
rect 283 -2105 330 -2071
rect 364 -2105 370 -2071
rect 162 -2143 370 -2105
rect 162 -2177 168 -2143
rect 202 -2177 249 -2143
rect 283 -2177 330 -2143
rect 364 -2177 370 -2143
rect 162 -2215 370 -2177
rect 162 -2249 168 -2215
rect 202 -2249 249 -2215
rect 283 -2249 330 -2215
rect 364 -2249 370 -2215
rect 162 -2287 370 -2249
rect 162 -2321 168 -2287
rect 202 -2321 249 -2287
rect 283 -2321 330 -2287
rect 364 -2321 370 -2287
rect 162 -2359 370 -2321
rect 162 -2393 168 -2359
rect 202 -2393 249 -2359
rect 283 -2393 330 -2359
rect 364 -2393 370 -2359
rect 162 -2431 370 -2393
rect 162 -2465 168 -2431
rect 202 -2465 249 -2431
rect 283 -2465 330 -2431
rect 364 -2465 370 -2431
rect 162 -2503 370 -2465
rect 162 -2537 168 -2503
rect 202 -2537 249 -2503
rect 283 -2537 330 -2503
rect 364 -2537 370 -2503
rect 162 -2575 370 -2537
rect 162 -2609 168 -2575
rect 202 -2609 249 -2575
rect 283 -2609 330 -2575
rect 364 -2609 370 -2575
rect 162 -2647 370 -2609
rect 162 -2681 168 -2647
rect 202 -2681 249 -2647
rect 283 -2681 330 -2647
rect 364 -2681 370 -2647
rect 162 -2719 370 -2681
rect 162 -2753 168 -2719
rect 202 -2753 249 -2719
rect 283 -2753 330 -2719
rect 364 -2753 370 -2719
rect 162 -2791 370 -2753
rect 162 -2825 168 -2791
rect 202 -2825 249 -2791
rect 283 -2825 330 -2791
rect 364 -2825 370 -2791
rect 162 -2863 370 -2825
rect 162 -2897 168 -2863
rect 202 -2897 249 -2863
rect 283 -2897 330 -2863
rect 364 -2897 370 -2863
rect 162 -2935 370 -2897
rect 162 -2969 168 -2935
rect 202 -2969 249 -2935
rect 283 -2969 330 -2935
rect 364 -2969 370 -2935
rect 162 -3007 370 -2969
rect 162 -3041 168 -3007
rect 202 -3041 249 -3007
rect 283 -3041 330 -3007
rect 364 -3041 370 -3007
rect 162 -3079 370 -3041
rect 162 -3113 168 -3079
rect 202 -3113 249 -3079
rect 283 -3113 330 -3079
rect 364 -3113 370 -3079
rect 162 -3151 370 -3113
rect 162 -3185 168 -3151
rect 202 -3185 249 -3151
rect 283 -3185 330 -3151
rect 364 -3185 370 -3151
rect 162 -3223 370 -3185
rect 162 -3257 168 -3223
rect 202 -3257 249 -3223
rect 283 -3257 330 -3223
rect 364 -3257 370 -3223
rect 162 -3295 370 -3257
rect 162 -3329 168 -3295
rect 202 -3329 249 -3295
rect 283 -3329 330 -3295
rect 364 -3329 370 -3295
rect 162 -3367 370 -3329
rect 162 -3401 168 -3367
rect 202 -3401 249 -3367
rect 283 -3401 330 -3367
rect 364 -3401 370 -3367
rect 162 -3439 370 -3401
rect 162 -3473 168 -3439
rect 202 -3473 249 -3439
rect 283 -3473 330 -3439
rect 364 -3473 370 -3439
rect 162 -3511 370 -3473
rect 162 -3545 168 -3511
rect 202 -3545 249 -3511
rect 283 -3545 330 -3511
rect 364 -3545 370 -3511
rect 162 -3583 370 -3545
rect 162 -3617 168 -3583
rect 202 -3617 249 -3583
rect 283 -3617 330 -3583
rect 364 -3617 370 -3583
rect 162 -3655 370 -3617
rect 162 -3689 168 -3655
rect 202 -3689 249 -3655
rect 283 -3689 330 -3655
rect 364 -3689 370 -3655
rect 162 -3727 370 -3689
rect 162 -3761 168 -3727
rect 202 -3761 249 -3727
rect 283 -3761 330 -3727
rect 364 -3761 370 -3727
rect 162 -3799 370 -3761
rect 162 -3833 168 -3799
rect 202 -3833 249 -3799
rect 283 -3833 330 -3799
rect 364 -3833 370 -3799
rect 162 -3871 370 -3833
rect 162 -3905 168 -3871
rect 202 -3905 249 -3871
rect 283 -3905 330 -3871
rect 364 -3905 370 -3871
rect 162 -3943 370 -3905
rect 162 -3977 168 -3943
rect 202 -3977 249 -3943
rect 283 -3977 330 -3943
rect 364 -3977 370 -3943
rect 162 -4015 370 -3977
rect 162 -4049 168 -4015
rect 202 -4049 249 -4015
rect 283 -4049 330 -4015
rect 364 -4049 370 -4015
rect 162 -4087 370 -4049
rect 162 -4121 168 -4087
rect 202 -4121 249 -4087
rect 283 -4121 330 -4087
rect 364 -4121 370 -4087
rect 162 -4159 370 -4121
rect 162 -4193 168 -4159
rect 202 -4193 249 -4159
rect 283 -4193 330 -4159
rect 364 -4193 370 -4159
rect 162 -4231 370 -4193
rect 162 -4265 168 -4231
rect 202 -4265 249 -4231
rect 283 -4265 330 -4231
rect 364 -4265 370 -4231
rect 162 -4303 370 -4265
rect 162 -4337 168 -4303
rect 202 -4337 249 -4303
rect 283 -4337 330 -4303
rect 364 -4337 370 -4303
rect 162 -4375 370 -4337
rect 162 -4409 168 -4375
rect 202 -4409 249 -4375
rect 283 -4409 330 -4375
rect 364 -4409 370 -4375
rect 162 -4447 370 -4409
rect 162 -4481 168 -4447
rect 202 -4481 249 -4447
rect 283 -4481 330 -4447
rect 364 -4481 370 -4447
rect 162 -4519 370 -4481
rect 162 -4553 168 -4519
rect 202 -4553 249 -4519
rect 283 -4553 330 -4519
rect 364 -4553 370 -4519
rect 162 -4591 370 -4553
rect 162 -4625 168 -4591
rect 202 -4625 249 -4591
rect 283 -4625 330 -4591
rect 364 -4625 370 -4591
rect 162 -4663 370 -4625
rect 162 -4697 168 -4663
rect 202 -4697 249 -4663
rect 283 -4697 330 -4663
rect 364 -4697 370 -4663
rect 162 -4735 370 -4697
rect 162 -4769 168 -4735
rect 202 -4769 249 -4735
rect 283 -4769 330 -4735
rect 364 -4769 370 -4735
rect 162 -4807 370 -4769
rect 162 -4841 168 -4807
rect 202 -4841 249 -4807
rect 283 -4841 330 -4807
rect 364 -4841 370 -4807
rect 162 -4879 370 -4841
rect 162 -4913 168 -4879
rect 202 -4913 249 -4879
rect 283 -4913 330 -4879
rect 364 -4913 370 -4879
rect 162 -4951 370 -4913
rect 162 -4985 168 -4951
rect 202 -4985 249 -4951
rect 283 -4985 330 -4951
rect 364 -4985 370 -4951
tri -162 -5062 -122 -5022 sw
tri 122 -5062 162 -5022 se
rect 162 -5062 370 -4985
tri 438 5000 458 5020 se
rect 458 5000 606 5020
tri 606 5000 626 5020 sw
rect 438 4985 626 5000
rect 438 -4985 479 4985
rect 585 -4985 626 4985
rect 438 -5000 626 -4985
tri 438 -5020 458 -5000 ne
rect 458 -5020 606 -5000
tri 606 -5020 626 -5000 nw
rect 694 4985 902 5062
tri 902 5022 942 5062 nw
tri 1186 5022 1226 5062 ne
rect 694 4951 700 4985
rect 734 4951 781 4985
rect 815 4951 862 4985
rect 896 4951 902 4985
rect 694 4913 902 4951
rect 694 4879 700 4913
rect 734 4879 781 4913
rect 815 4879 862 4913
rect 896 4879 902 4913
rect 694 4841 902 4879
rect 694 4807 700 4841
rect 734 4807 781 4841
rect 815 4807 862 4841
rect 896 4807 902 4841
rect 694 4769 902 4807
rect 694 4735 700 4769
rect 734 4735 781 4769
rect 815 4735 862 4769
rect 896 4735 902 4769
rect 694 4697 902 4735
rect 694 4663 700 4697
rect 734 4663 781 4697
rect 815 4663 862 4697
rect 896 4663 902 4697
rect 694 4625 902 4663
rect 694 4591 700 4625
rect 734 4591 781 4625
rect 815 4591 862 4625
rect 896 4591 902 4625
rect 694 4553 902 4591
rect 694 4519 700 4553
rect 734 4519 781 4553
rect 815 4519 862 4553
rect 896 4519 902 4553
rect 694 4481 902 4519
rect 694 4447 700 4481
rect 734 4447 781 4481
rect 815 4447 862 4481
rect 896 4447 902 4481
rect 694 4409 902 4447
rect 694 4375 700 4409
rect 734 4375 781 4409
rect 815 4375 862 4409
rect 896 4375 902 4409
rect 694 4337 902 4375
rect 694 4303 700 4337
rect 734 4303 781 4337
rect 815 4303 862 4337
rect 896 4303 902 4337
rect 694 4265 902 4303
rect 694 4231 700 4265
rect 734 4231 781 4265
rect 815 4231 862 4265
rect 896 4231 902 4265
rect 694 4193 902 4231
rect 694 4159 700 4193
rect 734 4159 781 4193
rect 815 4159 862 4193
rect 896 4159 902 4193
rect 694 4121 902 4159
rect 694 4087 700 4121
rect 734 4087 781 4121
rect 815 4087 862 4121
rect 896 4087 902 4121
rect 694 4049 902 4087
rect 694 4015 700 4049
rect 734 4015 781 4049
rect 815 4015 862 4049
rect 896 4015 902 4049
rect 694 3977 902 4015
rect 694 3943 700 3977
rect 734 3943 781 3977
rect 815 3943 862 3977
rect 896 3943 902 3977
rect 694 3905 902 3943
rect 694 3871 700 3905
rect 734 3871 781 3905
rect 815 3871 862 3905
rect 896 3871 902 3905
rect 694 3833 902 3871
rect 694 3799 700 3833
rect 734 3799 781 3833
rect 815 3799 862 3833
rect 896 3799 902 3833
rect 694 3761 902 3799
rect 694 3727 700 3761
rect 734 3727 781 3761
rect 815 3727 862 3761
rect 896 3727 902 3761
rect 694 3689 902 3727
rect 694 3655 700 3689
rect 734 3655 781 3689
rect 815 3655 862 3689
rect 896 3655 902 3689
rect 694 3617 902 3655
rect 694 3583 700 3617
rect 734 3583 781 3617
rect 815 3583 862 3617
rect 896 3583 902 3617
rect 694 3545 902 3583
rect 694 3511 700 3545
rect 734 3511 781 3545
rect 815 3511 862 3545
rect 896 3511 902 3545
rect 694 3473 902 3511
rect 694 3439 700 3473
rect 734 3439 781 3473
rect 815 3439 862 3473
rect 896 3439 902 3473
rect 694 3401 902 3439
rect 694 3367 700 3401
rect 734 3367 781 3401
rect 815 3367 862 3401
rect 896 3367 902 3401
rect 694 3329 902 3367
rect 694 3295 700 3329
rect 734 3295 781 3329
rect 815 3295 862 3329
rect 896 3295 902 3329
rect 694 3257 902 3295
rect 694 3223 700 3257
rect 734 3223 781 3257
rect 815 3223 862 3257
rect 896 3223 902 3257
rect 694 3185 902 3223
rect 694 3151 700 3185
rect 734 3151 781 3185
rect 815 3151 862 3185
rect 896 3151 902 3185
rect 694 3113 902 3151
rect 694 3079 700 3113
rect 734 3079 781 3113
rect 815 3079 862 3113
rect 896 3079 902 3113
rect 694 3041 902 3079
rect 694 3007 700 3041
rect 734 3007 781 3041
rect 815 3007 862 3041
rect 896 3007 902 3041
rect 694 2969 902 3007
rect 694 2935 700 2969
rect 734 2935 781 2969
rect 815 2935 862 2969
rect 896 2935 902 2969
rect 694 2897 902 2935
rect 694 2863 700 2897
rect 734 2863 781 2897
rect 815 2863 862 2897
rect 896 2863 902 2897
rect 694 2825 902 2863
rect 694 2791 700 2825
rect 734 2791 781 2825
rect 815 2791 862 2825
rect 896 2791 902 2825
rect 694 2753 902 2791
rect 694 2719 700 2753
rect 734 2719 781 2753
rect 815 2719 862 2753
rect 896 2719 902 2753
rect 694 2681 902 2719
rect 694 2647 700 2681
rect 734 2647 781 2681
rect 815 2647 862 2681
rect 896 2647 902 2681
rect 694 2609 902 2647
rect 694 2575 700 2609
rect 734 2575 781 2609
rect 815 2575 862 2609
rect 896 2575 902 2609
rect 694 2537 902 2575
rect 694 2503 700 2537
rect 734 2503 781 2537
rect 815 2503 862 2537
rect 896 2503 902 2537
rect 694 2465 902 2503
rect 694 2431 700 2465
rect 734 2431 781 2465
rect 815 2431 862 2465
rect 896 2431 902 2465
rect 694 2393 902 2431
rect 694 2359 700 2393
rect 734 2359 781 2393
rect 815 2359 862 2393
rect 896 2359 902 2393
rect 694 2321 902 2359
rect 694 2287 700 2321
rect 734 2287 781 2321
rect 815 2287 862 2321
rect 896 2287 902 2321
rect 694 2249 902 2287
rect 694 2215 700 2249
rect 734 2215 781 2249
rect 815 2215 862 2249
rect 896 2215 902 2249
rect 694 2177 902 2215
rect 694 2143 700 2177
rect 734 2143 781 2177
rect 815 2143 862 2177
rect 896 2143 902 2177
rect 694 2105 902 2143
rect 694 2071 700 2105
rect 734 2071 781 2105
rect 815 2071 862 2105
rect 896 2071 902 2105
rect 694 2033 902 2071
rect 694 1999 700 2033
rect 734 1999 781 2033
rect 815 1999 862 2033
rect 896 1999 902 2033
rect 694 1961 902 1999
rect 694 1927 700 1961
rect 734 1927 781 1961
rect 815 1927 862 1961
rect 896 1927 902 1961
rect 694 1889 902 1927
rect 694 1855 700 1889
rect 734 1855 781 1889
rect 815 1855 862 1889
rect 896 1855 902 1889
rect 694 1817 902 1855
rect 694 1783 700 1817
rect 734 1783 781 1817
rect 815 1783 862 1817
rect 896 1783 902 1817
rect 694 1745 902 1783
rect 694 1711 700 1745
rect 734 1711 781 1745
rect 815 1711 862 1745
rect 896 1711 902 1745
rect 694 1673 902 1711
rect 694 1639 700 1673
rect 734 1639 781 1673
rect 815 1639 862 1673
rect 896 1639 902 1673
rect 694 1601 902 1639
rect 694 1567 700 1601
rect 734 1567 781 1601
rect 815 1567 862 1601
rect 896 1567 902 1601
rect 694 1529 902 1567
rect 694 1495 700 1529
rect 734 1495 781 1529
rect 815 1495 862 1529
rect 896 1495 902 1529
rect 694 1457 902 1495
rect 694 1423 700 1457
rect 734 1423 781 1457
rect 815 1423 862 1457
rect 896 1423 902 1457
rect 694 1385 902 1423
rect 694 1351 700 1385
rect 734 1351 781 1385
rect 815 1351 862 1385
rect 896 1351 902 1385
rect 694 1313 902 1351
rect 694 1279 700 1313
rect 734 1279 781 1313
rect 815 1279 862 1313
rect 896 1279 902 1313
rect 694 1241 902 1279
rect 694 1207 700 1241
rect 734 1207 781 1241
rect 815 1207 862 1241
rect 896 1207 902 1241
rect 694 1169 902 1207
rect 694 1135 700 1169
rect 734 1135 781 1169
rect 815 1135 862 1169
rect 896 1135 902 1169
rect 694 1097 902 1135
rect 694 1063 700 1097
rect 734 1063 781 1097
rect 815 1063 862 1097
rect 896 1063 902 1097
rect 694 1025 902 1063
rect 694 991 700 1025
rect 734 991 781 1025
rect 815 991 862 1025
rect 896 991 902 1025
rect 694 953 902 991
rect 694 919 700 953
rect 734 919 781 953
rect 815 919 862 953
rect 896 919 902 953
rect 694 881 902 919
rect 694 847 700 881
rect 734 847 781 881
rect 815 847 862 881
rect 896 847 902 881
rect 694 809 902 847
rect 694 775 700 809
rect 734 775 781 809
rect 815 775 862 809
rect 896 775 902 809
rect 694 737 902 775
rect 694 703 700 737
rect 734 703 781 737
rect 815 703 862 737
rect 896 703 902 737
rect 694 665 902 703
rect 694 631 700 665
rect 734 631 781 665
rect 815 631 862 665
rect 896 631 902 665
rect 694 593 902 631
rect 694 559 700 593
rect 734 559 781 593
rect 815 559 862 593
rect 896 559 902 593
rect 694 521 902 559
rect 694 487 700 521
rect 734 487 781 521
rect 815 487 862 521
rect 896 487 902 521
rect 694 449 902 487
rect 694 415 700 449
rect 734 415 781 449
rect 815 415 862 449
rect 896 415 902 449
rect 694 377 902 415
rect 694 343 700 377
rect 734 343 781 377
rect 815 343 862 377
rect 896 343 902 377
rect 694 305 902 343
rect 694 271 700 305
rect 734 271 781 305
rect 815 271 862 305
rect 896 271 902 305
rect 694 233 902 271
rect 694 199 700 233
rect 734 199 781 233
rect 815 199 862 233
rect 896 199 902 233
rect 694 161 902 199
rect 694 127 700 161
rect 734 127 781 161
rect 815 127 862 161
rect 896 127 902 161
rect 694 89 902 127
rect 694 55 700 89
rect 734 55 781 89
rect 815 55 862 89
rect 896 55 902 89
rect 694 17 902 55
rect 694 -17 700 17
rect 734 -17 781 17
rect 815 -17 862 17
rect 896 -17 902 17
rect 694 -55 902 -17
rect 694 -89 700 -55
rect 734 -89 781 -55
rect 815 -89 862 -55
rect 896 -89 902 -55
rect 694 -127 902 -89
rect 694 -161 700 -127
rect 734 -161 781 -127
rect 815 -161 862 -127
rect 896 -161 902 -127
rect 694 -199 902 -161
rect 694 -233 700 -199
rect 734 -233 781 -199
rect 815 -233 862 -199
rect 896 -233 902 -199
rect 694 -271 902 -233
rect 694 -305 700 -271
rect 734 -305 781 -271
rect 815 -305 862 -271
rect 896 -305 902 -271
rect 694 -343 902 -305
rect 694 -377 700 -343
rect 734 -377 781 -343
rect 815 -377 862 -343
rect 896 -377 902 -343
rect 694 -415 902 -377
rect 694 -449 700 -415
rect 734 -449 781 -415
rect 815 -449 862 -415
rect 896 -449 902 -415
rect 694 -487 902 -449
rect 694 -521 700 -487
rect 734 -521 781 -487
rect 815 -521 862 -487
rect 896 -521 902 -487
rect 694 -559 902 -521
rect 694 -593 700 -559
rect 734 -593 781 -559
rect 815 -593 862 -559
rect 896 -593 902 -559
rect 694 -631 902 -593
rect 694 -665 700 -631
rect 734 -665 781 -631
rect 815 -665 862 -631
rect 896 -665 902 -631
rect 694 -703 902 -665
rect 694 -737 700 -703
rect 734 -737 781 -703
rect 815 -737 862 -703
rect 896 -737 902 -703
rect 694 -775 902 -737
rect 694 -809 700 -775
rect 734 -809 781 -775
rect 815 -809 862 -775
rect 896 -809 902 -775
rect 694 -847 902 -809
rect 694 -881 700 -847
rect 734 -881 781 -847
rect 815 -881 862 -847
rect 896 -881 902 -847
rect 694 -919 902 -881
rect 694 -953 700 -919
rect 734 -953 781 -919
rect 815 -953 862 -919
rect 896 -953 902 -919
rect 694 -991 902 -953
rect 694 -1025 700 -991
rect 734 -1025 781 -991
rect 815 -1025 862 -991
rect 896 -1025 902 -991
rect 694 -1063 902 -1025
rect 694 -1097 700 -1063
rect 734 -1097 781 -1063
rect 815 -1097 862 -1063
rect 896 -1097 902 -1063
rect 694 -1135 902 -1097
rect 694 -1169 700 -1135
rect 734 -1169 781 -1135
rect 815 -1169 862 -1135
rect 896 -1169 902 -1135
rect 694 -1207 902 -1169
rect 694 -1241 700 -1207
rect 734 -1241 781 -1207
rect 815 -1241 862 -1207
rect 896 -1241 902 -1207
rect 694 -1279 902 -1241
rect 694 -1313 700 -1279
rect 734 -1313 781 -1279
rect 815 -1313 862 -1279
rect 896 -1313 902 -1279
rect 694 -1351 902 -1313
rect 694 -1385 700 -1351
rect 734 -1385 781 -1351
rect 815 -1385 862 -1351
rect 896 -1385 902 -1351
rect 694 -1423 902 -1385
rect 694 -1457 700 -1423
rect 734 -1457 781 -1423
rect 815 -1457 862 -1423
rect 896 -1457 902 -1423
rect 694 -1495 902 -1457
rect 694 -1529 700 -1495
rect 734 -1529 781 -1495
rect 815 -1529 862 -1495
rect 896 -1529 902 -1495
rect 694 -1567 902 -1529
rect 694 -1601 700 -1567
rect 734 -1601 781 -1567
rect 815 -1601 862 -1567
rect 896 -1601 902 -1567
rect 694 -1639 902 -1601
rect 694 -1673 700 -1639
rect 734 -1673 781 -1639
rect 815 -1673 862 -1639
rect 896 -1673 902 -1639
rect 694 -1711 902 -1673
rect 694 -1745 700 -1711
rect 734 -1745 781 -1711
rect 815 -1745 862 -1711
rect 896 -1745 902 -1711
rect 694 -1783 902 -1745
rect 694 -1817 700 -1783
rect 734 -1817 781 -1783
rect 815 -1817 862 -1783
rect 896 -1817 902 -1783
rect 694 -1855 902 -1817
rect 694 -1889 700 -1855
rect 734 -1889 781 -1855
rect 815 -1889 862 -1855
rect 896 -1889 902 -1855
rect 694 -1927 902 -1889
rect 694 -1961 700 -1927
rect 734 -1961 781 -1927
rect 815 -1961 862 -1927
rect 896 -1961 902 -1927
rect 694 -1999 902 -1961
rect 694 -2033 700 -1999
rect 734 -2033 781 -1999
rect 815 -2033 862 -1999
rect 896 -2033 902 -1999
rect 694 -2071 902 -2033
rect 694 -2105 700 -2071
rect 734 -2105 781 -2071
rect 815 -2105 862 -2071
rect 896 -2105 902 -2071
rect 694 -2143 902 -2105
rect 694 -2177 700 -2143
rect 734 -2177 781 -2143
rect 815 -2177 862 -2143
rect 896 -2177 902 -2143
rect 694 -2215 902 -2177
rect 694 -2249 700 -2215
rect 734 -2249 781 -2215
rect 815 -2249 862 -2215
rect 896 -2249 902 -2215
rect 694 -2287 902 -2249
rect 694 -2321 700 -2287
rect 734 -2321 781 -2287
rect 815 -2321 862 -2287
rect 896 -2321 902 -2287
rect 694 -2359 902 -2321
rect 694 -2393 700 -2359
rect 734 -2393 781 -2359
rect 815 -2393 862 -2359
rect 896 -2393 902 -2359
rect 694 -2431 902 -2393
rect 694 -2465 700 -2431
rect 734 -2465 781 -2431
rect 815 -2465 862 -2431
rect 896 -2465 902 -2431
rect 694 -2503 902 -2465
rect 694 -2537 700 -2503
rect 734 -2537 781 -2503
rect 815 -2537 862 -2503
rect 896 -2537 902 -2503
rect 694 -2575 902 -2537
rect 694 -2609 700 -2575
rect 734 -2609 781 -2575
rect 815 -2609 862 -2575
rect 896 -2609 902 -2575
rect 694 -2647 902 -2609
rect 694 -2681 700 -2647
rect 734 -2681 781 -2647
rect 815 -2681 862 -2647
rect 896 -2681 902 -2647
rect 694 -2719 902 -2681
rect 694 -2753 700 -2719
rect 734 -2753 781 -2719
rect 815 -2753 862 -2719
rect 896 -2753 902 -2719
rect 694 -2791 902 -2753
rect 694 -2825 700 -2791
rect 734 -2825 781 -2791
rect 815 -2825 862 -2791
rect 896 -2825 902 -2791
rect 694 -2863 902 -2825
rect 694 -2897 700 -2863
rect 734 -2897 781 -2863
rect 815 -2897 862 -2863
rect 896 -2897 902 -2863
rect 694 -2935 902 -2897
rect 694 -2969 700 -2935
rect 734 -2969 781 -2935
rect 815 -2969 862 -2935
rect 896 -2969 902 -2935
rect 694 -3007 902 -2969
rect 694 -3041 700 -3007
rect 734 -3041 781 -3007
rect 815 -3041 862 -3007
rect 896 -3041 902 -3007
rect 694 -3079 902 -3041
rect 694 -3113 700 -3079
rect 734 -3113 781 -3079
rect 815 -3113 862 -3079
rect 896 -3113 902 -3079
rect 694 -3151 902 -3113
rect 694 -3185 700 -3151
rect 734 -3185 781 -3151
rect 815 -3185 862 -3151
rect 896 -3185 902 -3151
rect 694 -3223 902 -3185
rect 694 -3257 700 -3223
rect 734 -3257 781 -3223
rect 815 -3257 862 -3223
rect 896 -3257 902 -3223
rect 694 -3295 902 -3257
rect 694 -3329 700 -3295
rect 734 -3329 781 -3295
rect 815 -3329 862 -3295
rect 896 -3329 902 -3295
rect 694 -3367 902 -3329
rect 694 -3401 700 -3367
rect 734 -3401 781 -3367
rect 815 -3401 862 -3367
rect 896 -3401 902 -3367
rect 694 -3439 902 -3401
rect 694 -3473 700 -3439
rect 734 -3473 781 -3439
rect 815 -3473 862 -3439
rect 896 -3473 902 -3439
rect 694 -3511 902 -3473
rect 694 -3545 700 -3511
rect 734 -3545 781 -3511
rect 815 -3545 862 -3511
rect 896 -3545 902 -3511
rect 694 -3583 902 -3545
rect 694 -3617 700 -3583
rect 734 -3617 781 -3583
rect 815 -3617 862 -3583
rect 896 -3617 902 -3583
rect 694 -3655 902 -3617
rect 694 -3689 700 -3655
rect 734 -3689 781 -3655
rect 815 -3689 862 -3655
rect 896 -3689 902 -3655
rect 694 -3727 902 -3689
rect 694 -3761 700 -3727
rect 734 -3761 781 -3727
rect 815 -3761 862 -3727
rect 896 -3761 902 -3727
rect 694 -3799 902 -3761
rect 694 -3833 700 -3799
rect 734 -3833 781 -3799
rect 815 -3833 862 -3799
rect 896 -3833 902 -3799
rect 694 -3871 902 -3833
rect 694 -3905 700 -3871
rect 734 -3905 781 -3871
rect 815 -3905 862 -3871
rect 896 -3905 902 -3871
rect 694 -3943 902 -3905
rect 694 -3977 700 -3943
rect 734 -3977 781 -3943
rect 815 -3977 862 -3943
rect 896 -3977 902 -3943
rect 694 -4015 902 -3977
rect 694 -4049 700 -4015
rect 734 -4049 781 -4015
rect 815 -4049 862 -4015
rect 896 -4049 902 -4015
rect 694 -4087 902 -4049
rect 694 -4121 700 -4087
rect 734 -4121 781 -4087
rect 815 -4121 862 -4087
rect 896 -4121 902 -4087
rect 694 -4159 902 -4121
rect 694 -4193 700 -4159
rect 734 -4193 781 -4159
rect 815 -4193 862 -4159
rect 896 -4193 902 -4159
rect 694 -4231 902 -4193
rect 694 -4265 700 -4231
rect 734 -4265 781 -4231
rect 815 -4265 862 -4231
rect 896 -4265 902 -4231
rect 694 -4303 902 -4265
rect 694 -4337 700 -4303
rect 734 -4337 781 -4303
rect 815 -4337 862 -4303
rect 896 -4337 902 -4303
rect 694 -4375 902 -4337
rect 694 -4409 700 -4375
rect 734 -4409 781 -4375
rect 815 -4409 862 -4375
rect 896 -4409 902 -4375
rect 694 -4447 902 -4409
rect 694 -4481 700 -4447
rect 734 -4481 781 -4447
rect 815 -4481 862 -4447
rect 896 -4481 902 -4447
rect 694 -4519 902 -4481
rect 694 -4553 700 -4519
rect 734 -4553 781 -4519
rect 815 -4553 862 -4519
rect 896 -4553 902 -4519
rect 694 -4591 902 -4553
rect 694 -4625 700 -4591
rect 734 -4625 781 -4591
rect 815 -4625 862 -4591
rect 896 -4625 902 -4591
rect 694 -4663 902 -4625
rect 694 -4697 700 -4663
rect 734 -4697 781 -4663
rect 815 -4697 862 -4663
rect 896 -4697 902 -4663
rect 694 -4735 902 -4697
rect 694 -4769 700 -4735
rect 734 -4769 781 -4735
rect 815 -4769 862 -4735
rect 896 -4769 902 -4735
rect 694 -4807 902 -4769
rect 694 -4841 700 -4807
rect 734 -4841 781 -4807
rect 815 -4841 862 -4807
rect 896 -4841 902 -4807
rect 694 -4879 902 -4841
rect 694 -4913 700 -4879
rect 734 -4913 781 -4879
rect 815 -4913 862 -4879
rect 896 -4913 902 -4879
rect 694 -4951 902 -4913
rect 694 -4985 700 -4951
rect 734 -4985 781 -4951
rect 815 -4985 862 -4951
rect 896 -4985 902 -4951
tri 370 -5062 410 -5022 sw
tri 654 -5062 694 -5022 se
rect 694 -5062 902 -4985
tri 970 5000 990 5020 se
rect 990 5000 1138 5020
tri 1138 5000 1158 5020 sw
rect 970 4985 1158 5000
rect 970 -4985 1011 4985
rect 1117 -4985 1158 4985
rect 970 -5000 1158 -4985
tri 970 -5020 990 -5000 ne
rect 990 -5020 1138 -5000
tri 1138 -5020 1158 -5000 nw
rect 1226 4985 1330 5062
rect 1226 4951 1232 4985
rect 1266 4951 1330 4985
rect 1226 4913 1330 4951
rect 1226 4879 1232 4913
rect 1266 4879 1330 4913
rect 1226 4841 1330 4879
rect 1226 4807 1232 4841
rect 1266 4807 1330 4841
rect 1226 4769 1330 4807
rect 1226 4735 1232 4769
rect 1266 4735 1330 4769
rect 1226 4697 1330 4735
rect 1226 4663 1232 4697
rect 1266 4663 1330 4697
rect 1226 4625 1330 4663
rect 1226 4591 1232 4625
rect 1266 4591 1330 4625
rect 1226 4553 1330 4591
rect 1226 4519 1232 4553
rect 1266 4519 1330 4553
rect 1226 4481 1330 4519
rect 1226 4447 1232 4481
rect 1266 4447 1330 4481
rect 1226 4409 1330 4447
rect 1226 4375 1232 4409
rect 1266 4375 1330 4409
rect 1226 4337 1330 4375
rect 1226 4303 1232 4337
rect 1266 4303 1330 4337
rect 1226 4265 1330 4303
rect 1226 4231 1232 4265
rect 1266 4231 1330 4265
rect 1226 4193 1330 4231
rect 1226 4159 1232 4193
rect 1266 4159 1330 4193
rect 1226 4121 1330 4159
rect 1226 4087 1232 4121
rect 1266 4087 1330 4121
rect 1226 4049 1330 4087
rect 1226 4015 1232 4049
rect 1266 4015 1330 4049
rect 1226 3977 1330 4015
rect 1226 3943 1232 3977
rect 1266 3943 1330 3977
rect 1226 3905 1330 3943
rect 1226 3871 1232 3905
rect 1266 3871 1330 3905
rect 1226 3833 1330 3871
rect 1226 3799 1232 3833
rect 1266 3799 1330 3833
rect 1226 3761 1330 3799
rect 1226 3727 1232 3761
rect 1266 3727 1330 3761
rect 1226 3689 1330 3727
rect 1226 3655 1232 3689
rect 1266 3655 1330 3689
rect 1226 3617 1330 3655
rect 1226 3583 1232 3617
rect 1266 3583 1330 3617
rect 1226 3545 1330 3583
rect 1226 3511 1232 3545
rect 1266 3511 1330 3545
rect 1226 3473 1330 3511
rect 1226 3439 1232 3473
rect 1266 3439 1330 3473
rect 1226 3401 1330 3439
rect 1226 3367 1232 3401
rect 1266 3367 1330 3401
rect 1226 3329 1330 3367
rect 1226 3295 1232 3329
rect 1266 3295 1330 3329
rect 1226 3257 1330 3295
rect 1226 3223 1232 3257
rect 1266 3223 1330 3257
rect 1226 3185 1330 3223
rect 1226 3151 1232 3185
rect 1266 3151 1330 3185
rect 1226 3113 1330 3151
rect 1226 3079 1232 3113
rect 1266 3079 1330 3113
rect 1226 3041 1330 3079
rect 1226 3007 1232 3041
rect 1266 3007 1330 3041
rect 1226 2969 1330 3007
rect 1226 2935 1232 2969
rect 1266 2935 1330 2969
rect 1226 2897 1330 2935
rect 1226 2863 1232 2897
rect 1266 2863 1330 2897
rect 1226 2825 1330 2863
rect 1226 2791 1232 2825
rect 1266 2791 1330 2825
rect 1226 2753 1330 2791
rect 1226 2719 1232 2753
rect 1266 2719 1330 2753
rect 1226 2681 1330 2719
rect 1226 2647 1232 2681
rect 1266 2647 1330 2681
rect 1226 2609 1330 2647
rect 1226 2575 1232 2609
rect 1266 2575 1330 2609
rect 1226 2537 1330 2575
rect 1226 2503 1232 2537
rect 1266 2503 1330 2537
rect 1226 2465 1330 2503
rect 1226 2431 1232 2465
rect 1266 2431 1330 2465
rect 1226 2393 1330 2431
rect 1226 2359 1232 2393
rect 1266 2359 1330 2393
rect 1226 2321 1330 2359
rect 1226 2287 1232 2321
rect 1266 2287 1330 2321
rect 1226 2249 1330 2287
rect 1226 2215 1232 2249
rect 1266 2215 1330 2249
rect 1226 2177 1330 2215
rect 1226 2143 1232 2177
rect 1266 2143 1330 2177
rect 1226 2105 1330 2143
rect 1226 2071 1232 2105
rect 1266 2071 1330 2105
rect 1226 2033 1330 2071
rect 1226 1999 1232 2033
rect 1266 1999 1330 2033
rect 1226 1961 1330 1999
rect 1226 1927 1232 1961
rect 1266 1927 1330 1961
rect 1226 1889 1330 1927
rect 1226 1855 1232 1889
rect 1266 1855 1330 1889
rect 1226 1817 1330 1855
rect 1226 1783 1232 1817
rect 1266 1783 1330 1817
rect 1226 1745 1330 1783
rect 1226 1711 1232 1745
rect 1266 1711 1330 1745
rect 1226 1673 1330 1711
rect 1226 1639 1232 1673
rect 1266 1639 1330 1673
rect 1226 1601 1330 1639
rect 1226 1567 1232 1601
rect 1266 1567 1330 1601
rect 1226 1529 1330 1567
rect 1226 1495 1232 1529
rect 1266 1495 1330 1529
rect 1226 1457 1330 1495
rect 1226 1423 1232 1457
rect 1266 1423 1330 1457
rect 1226 1385 1330 1423
rect 1226 1351 1232 1385
rect 1266 1351 1330 1385
rect 1226 1313 1330 1351
rect 1226 1279 1232 1313
rect 1266 1279 1330 1313
rect 1226 1241 1330 1279
rect 1226 1207 1232 1241
rect 1266 1207 1330 1241
rect 1226 1169 1330 1207
rect 1226 1135 1232 1169
rect 1266 1135 1330 1169
rect 1226 1097 1330 1135
rect 1226 1063 1232 1097
rect 1266 1063 1330 1097
rect 1226 1025 1330 1063
rect 1226 991 1232 1025
rect 1266 991 1330 1025
rect 1226 953 1330 991
rect 1226 919 1232 953
rect 1266 919 1330 953
rect 1226 881 1330 919
rect 1226 847 1232 881
rect 1266 847 1330 881
rect 1226 809 1330 847
rect 1226 775 1232 809
rect 1266 775 1330 809
rect 1226 737 1330 775
rect 1226 703 1232 737
rect 1266 703 1330 737
rect 1226 665 1330 703
rect 1226 631 1232 665
rect 1266 631 1330 665
rect 1226 593 1330 631
rect 1226 559 1232 593
rect 1266 559 1330 593
rect 1226 521 1330 559
rect 1226 487 1232 521
rect 1266 487 1330 521
rect 1226 449 1330 487
rect 1226 415 1232 449
rect 1266 415 1330 449
rect 1226 377 1330 415
rect 1226 343 1232 377
rect 1266 343 1330 377
rect 1226 305 1330 343
rect 1226 271 1232 305
rect 1266 271 1330 305
rect 1226 233 1330 271
rect 1226 199 1232 233
rect 1266 199 1330 233
rect 1226 161 1330 199
rect 1226 127 1232 161
rect 1266 127 1330 161
rect 1226 89 1330 127
rect 1226 55 1232 89
rect 1266 55 1330 89
rect 1226 17 1330 55
rect 1226 -17 1232 17
rect 1266 -17 1330 17
rect 1226 -55 1330 -17
rect 1226 -89 1232 -55
rect 1266 -89 1330 -55
rect 1226 -127 1330 -89
rect 1226 -161 1232 -127
rect 1266 -161 1330 -127
rect 1226 -199 1330 -161
rect 1226 -233 1232 -199
rect 1266 -233 1330 -199
rect 1226 -271 1330 -233
rect 1226 -305 1232 -271
rect 1266 -305 1330 -271
rect 1226 -343 1330 -305
rect 1226 -377 1232 -343
rect 1266 -377 1330 -343
rect 1226 -415 1330 -377
rect 1226 -449 1232 -415
rect 1266 -449 1330 -415
rect 1226 -487 1330 -449
rect 1226 -521 1232 -487
rect 1266 -521 1330 -487
rect 1226 -559 1330 -521
rect 1226 -593 1232 -559
rect 1266 -593 1330 -559
rect 1226 -631 1330 -593
rect 1226 -665 1232 -631
rect 1266 -665 1330 -631
rect 1226 -703 1330 -665
rect 1226 -737 1232 -703
rect 1266 -737 1330 -703
rect 1226 -775 1330 -737
rect 1226 -809 1232 -775
rect 1266 -809 1330 -775
rect 1226 -847 1330 -809
rect 1226 -881 1232 -847
rect 1266 -881 1330 -847
rect 1226 -919 1330 -881
rect 1226 -953 1232 -919
rect 1266 -953 1330 -919
rect 1226 -991 1330 -953
rect 1226 -1025 1232 -991
rect 1266 -1025 1330 -991
rect 1226 -1063 1330 -1025
rect 1226 -1097 1232 -1063
rect 1266 -1097 1330 -1063
rect 1226 -1135 1330 -1097
rect 1226 -1169 1232 -1135
rect 1266 -1169 1330 -1135
rect 1226 -1207 1330 -1169
rect 1226 -1241 1232 -1207
rect 1266 -1241 1330 -1207
rect 1226 -1279 1330 -1241
rect 1226 -1313 1232 -1279
rect 1266 -1313 1330 -1279
rect 1226 -1351 1330 -1313
rect 1226 -1385 1232 -1351
rect 1266 -1385 1330 -1351
rect 1226 -1423 1330 -1385
rect 1226 -1457 1232 -1423
rect 1266 -1457 1330 -1423
rect 1226 -1495 1330 -1457
rect 1226 -1529 1232 -1495
rect 1266 -1529 1330 -1495
rect 1226 -1567 1330 -1529
rect 1226 -1601 1232 -1567
rect 1266 -1601 1330 -1567
rect 1226 -1639 1330 -1601
rect 1226 -1673 1232 -1639
rect 1266 -1673 1330 -1639
rect 1226 -1711 1330 -1673
rect 1226 -1745 1232 -1711
rect 1266 -1745 1330 -1711
rect 1226 -1783 1330 -1745
rect 1226 -1817 1232 -1783
rect 1266 -1817 1330 -1783
rect 1226 -1855 1330 -1817
rect 1226 -1889 1232 -1855
rect 1266 -1889 1330 -1855
rect 1226 -1927 1330 -1889
rect 1226 -1961 1232 -1927
rect 1266 -1961 1330 -1927
rect 1226 -1999 1330 -1961
rect 1226 -2033 1232 -1999
rect 1266 -2033 1330 -1999
rect 1226 -2071 1330 -2033
rect 1226 -2105 1232 -2071
rect 1266 -2105 1330 -2071
rect 1226 -2143 1330 -2105
rect 1226 -2177 1232 -2143
rect 1266 -2177 1330 -2143
rect 1226 -2215 1330 -2177
rect 1226 -2249 1232 -2215
rect 1266 -2249 1330 -2215
rect 1226 -2287 1330 -2249
rect 1226 -2321 1232 -2287
rect 1266 -2321 1330 -2287
rect 1226 -2359 1330 -2321
rect 1226 -2393 1232 -2359
rect 1266 -2393 1330 -2359
rect 1226 -2431 1330 -2393
rect 1226 -2465 1232 -2431
rect 1266 -2465 1330 -2431
rect 1226 -2503 1330 -2465
rect 1226 -2537 1232 -2503
rect 1266 -2537 1330 -2503
rect 1226 -2575 1330 -2537
rect 1226 -2609 1232 -2575
rect 1266 -2609 1330 -2575
rect 1226 -2647 1330 -2609
rect 1226 -2681 1232 -2647
rect 1266 -2681 1330 -2647
rect 1226 -2719 1330 -2681
rect 1226 -2753 1232 -2719
rect 1266 -2753 1330 -2719
rect 1226 -2791 1330 -2753
rect 1226 -2825 1232 -2791
rect 1266 -2825 1330 -2791
rect 1226 -2863 1330 -2825
rect 1226 -2897 1232 -2863
rect 1266 -2897 1330 -2863
rect 1226 -2935 1330 -2897
rect 1226 -2969 1232 -2935
rect 1266 -2969 1330 -2935
rect 1226 -3007 1330 -2969
rect 1226 -3041 1232 -3007
rect 1266 -3041 1330 -3007
rect 1226 -3079 1330 -3041
rect 1226 -3113 1232 -3079
rect 1266 -3113 1330 -3079
rect 1226 -3151 1330 -3113
rect 1226 -3185 1232 -3151
rect 1266 -3185 1330 -3151
rect 1226 -3223 1330 -3185
rect 1226 -3257 1232 -3223
rect 1266 -3257 1330 -3223
rect 1226 -3295 1330 -3257
rect 1226 -3329 1232 -3295
rect 1266 -3329 1330 -3295
rect 1226 -3367 1330 -3329
rect 1226 -3401 1232 -3367
rect 1266 -3401 1330 -3367
rect 1226 -3439 1330 -3401
rect 1226 -3473 1232 -3439
rect 1266 -3473 1330 -3439
rect 1226 -3511 1330 -3473
rect 1226 -3545 1232 -3511
rect 1266 -3545 1330 -3511
rect 1226 -3583 1330 -3545
rect 1226 -3617 1232 -3583
rect 1266 -3617 1330 -3583
rect 1226 -3655 1330 -3617
rect 1226 -3689 1232 -3655
rect 1266 -3689 1330 -3655
rect 1226 -3727 1330 -3689
rect 1226 -3761 1232 -3727
rect 1266 -3761 1330 -3727
rect 1226 -3799 1330 -3761
rect 1226 -3833 1232 -3799
rect 1266 -3833 1330 -3799
rect 1226 -3871 1330 -3833
rect 1226 -3905 1232 -3871
rect 1266 -3905 1330 -3871
rect 1226 -3943 1330 -3905
rect 1226 -3977 1232 -3943
rect 1266 -3977 1330 -3943
rect 1226 -4015 1330 -3977
rect 1226 -4049 1232 -4015
rect 1266 -4049 1330 -4015
rect 1226 -4087 1330 -4049
rect 1226 -4121 1232 -4087
rect 1266 -4121 1330 -4087
rect 1226 -4159 1330 -4121
rect 1226 -4193 1232 -4159
rect 1266 -4193 1330 -4159
rect 1226 -4231 1330 -4193
rect 1226 -4265 1232 -4231
rect 1266 -4265 1330 -4231
rect 1226 -4303 1330 -4265
rect 1226 -4337 1232 -4303
rect 1266 -4337 1330 -4303
rect 1226 -4375 1330 -4337
rect 1226 -4409 1232 -4375
rect 1266 -4409 1330 -4375
rect 1226 -4447 1330 -4409
rect 1226 -4481 1232 -4447
rect 1266 -4481 1330 -4447
rect 1226 -4519 1330 -4481
rect 1226 -4553 1232 -4519
rect 1266 -4553 1330 -4519
rect 1226 -4591 1330 -4553
rect 1226 -4625 1232 -4591
rect 1266 -4625 1330 -4591
rect 1226 -4663 1330 -4625
rect 1226 -4697 1232 -4663
rect 1266 -4697 1330 -4663
rect 1226 -4735 1330 -4697
rect 1226 -4769 1232 -4735
rect 1266 -4769 1330 -4735
rect 1226 -4807 1330 -4769
rect 1226 -4841 1232 -4807
rect 1266 -4841 1330 -4807
rect 1226 -4879 1330 -4841
rect 1226 -4913 1232 -4879
rect 1266 -4913 1330 -4879
rect 1226 -4951 1330 -4913
rect 1226 -4985 1232 -4951
rect 1266 -4985 1330 -4951
tri 902 -5062 942 -5022 sw
tri 1186 -5062 1226 -5022 se
rect 1226 -5062 1330 -4985
rect -1330 -5068 1330 -5062
rect -1330 -5102 -1153 -5068
rect -1119 -5102 -1081 -5068
rect -1047 -5102 -1009 -5068
rect -975 -5102 -621 -5068
rect -587 -5102 -549 -5068
rect -515 -5102 -477 -5068
rect -443 -5102 -89 -5068
rect -55 -5102 -17 -5068
rect 17 -5102 55 -5068
rect 89 -5102 443 -5068
rect 477 -5102 515 -5068
rect 549 -5102 587 -5068
rect 621 -5102 975 -5068
rect 1009 -5102 1047 -5068
rect 1081 -5102 1119 -5068
rect 1153 -5102 1330 -5068
rect -1330 -5168 1330 -5102
rect -1956 -5268 -1493 -5237
rect 1488 -5237 1542 5237
rect 1936 -5237 1956 5237
tri -1493 -5268 -1471 -5246 sw
tri 1466 -5268 1488 -5246 se
rect 1488 -5268 1956 -5237
rect -1956 -5286 -1471 -5268
tri -1471 -5286 -1453 -5268 sw
tri 1448 -5286 1466 -5268 se
rect 1466 -5286 1956 -5268
rect -1956 -5346 1956 -5286
rect -1956 -5360 -1421 -5346
tri -1956 -5740 -1576 -5360 ne
rect -1576 -5740 -1421 -5360
rect 1421 -5360 1956 -5346
rect 1421 -5740 1556 -5360
tri -1576 -5760 -1556 -5740 ne
rect -1556 -5760 1556 -5740
tri 1556 -5760 1956 -5360 nw
<< properties >>
string FIXED_BBOX 879 -5085 1249 5085
string GDS_END 2376950
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__analog.gds
string GDS_START 1582434
<< end >>
