magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< obsli1 >>
rect 385 961 1913 980
rect 190 817 256 883
rect 385 855 412 961
rect 1886 855 1913 961
rect 385 843 1913 855
rect 2042 817 2108 883
rect 190 795 230 817
rect 2068 795 2108 817
rect 41 759 230 795
rect 41 725 60 759
rect 94 725 230 759
rect 41 687 230 725
rect 41 653 60 687
rect 94 653 230 687
rect 41 615 230 653
rect 41 581 60 615
rect 94 581 230 615
rect 41 543 230 581
rect 41 509 60 543
rect 94 509 230 543
rect 41 471 230 509
rect 41 437 60 471
rect 94 437 230 471
rect 41 399 230 437
rect 41 365 60 399
rect 94 365 230 399
rect 41 327 230 365
rect 41 293 60 327
rect 94 293 230 327
rect 41 255 230 293
rect 41 221 60 255
rect 94 221 230 255
rect 41 185 230 221
rect 352 185 386 795
rect 508 185 542 795
rect 664 185 698 795
rect 820 185 854 795
rect 976 185 1010 795
rect 1132 185 1166 795
rect 1288 185 1322 795
rect 1444 185 1478 795
rect 1600 185 1634 795
rect 1756 185 1790 795
rect 1912 185 1946 795
rect 2068 759 2257 795
rect 2068 725 2204 759
rect 2238 725 2257 759
rect 2068 687 2257 725
rect 2068 653 2204 687
rect 2238 653 2257 687
rect 2068 615 2257 653
rect 2068 581 2204 615
rect 2238 581 2257 615
rect 2068 543 2257 581
rect 2068 509 2204 543
rect 2238 509 2257 543
rect 2068 471 2257 509
rect 2068 437 2204 471
rect 2238 437 2257 471
rect 2068 399 2257 437
rect 2068 365 2204 399
rect 2238 365 2257 399
rect 2068 327 2257 365
rect 2068 293 2204 327
rect 2238 293 2257 327
rect 2068 255 2257 293
rect 2068 221 2204 255
rect 2238 221 2257 255
rect 2068 185 2257 221
rect 190 163 230 185
rect 2068 163 2108 185
rect 190 97 256 163
rect 385 125 1913 137
rect 385 19 412 125
rect 1886 19 1913 125
rect 2042 97 2108 163
rect 385 0 1913 19
<< obsli1c >>
rect 412 855 1886 961
rect 60 725 94 759
rect 60 653 94 687
rect 60 581 94 615
rect 60 509 94 543
rect 60 437 94 471
rect 60 365 94 399
rect 60 293 94 327
rect 60 221 94 255
rect 2204 725 2238 759
rect 2204 653 2238 687
rect 2204 581 2238 615
rect 2204 509 2238 543
rect 2204 437 2238 471
rect 2204 365 2238 399
rect 2204 293 2238 327
rect 2204 221 2238 255
rect 412 19 1886 125
<< metal1 >>
rect 381 961 1917 980
rect 381 855 412 961
rect 1886 855 1917 961
rect 381 843 1917 855
rect 41 759 100 771
rect 41 725 60 759
rect 94 725 100 759
rect 41 687 100 725
rect 41 653 60 687
rect 94 653 100 687
rect 41 615 100 653
rect 41 581 60 615
rect 94 581 100 615
rect 41 543 100 581
rect 41 509 60 543
rect 94 509 100 543
rect 41 471 100 509
rect 41 437 60 471
rect 94 437 100 471
rect 41 399 100 437
rect 41 365 60 399
rect 94 365 100 399
rect 41 327 100 365
rect 41 293 60 327
rect 94 293 100 327
rect 41 255 100 293
rect 41 221 60 255
rect 94 221 100 255
rect 41 209 100 221
rect 2198 759 2257 771
rect 2198 725 2204 759
rect 2238 725 2257 759
rect 2198 687 2257 725
rect 2198 653 2204 687
rect 2238 653 2257 687
rect 2198 615 2257 653
rect 2198 581 2204 615
rect 2238 581 2257 615
rect 2198 543 2257 581
rect 2198 509 2204 543
rect 2238 509 2257 543
rect 2198 471 2257 509
rect 2198 437 2204 471
rect 2238 437 2257 471
rect 2198 399 2257 437
rect 2198 365 2204 399
rect 2238 365 2257 399
rect 2198 327 2257 365
rect 2198 293 2204 327
rect 2238 293 2257 327
rect 2198 255 2257 293
rect 2198 221 2204 255
rect 2238 221 2257 255
rect 2198 209 2257 221
rect 381 125 1917 137
rect 381 19 412 125
rect 1886 19 1917 125
rect 381 0 1917 19
<< obsm1 >>
rect 343 209 395 771
rect 499 209 551 771
rect 655 209 707 771
rect 811 209 863 771
rect 967 209 1019 771
rect 1123 209 1175 771
rect 1279 209 1331 771
rect 1435 209 1487 771
rect 1591 209 1643 771
rect 1747 209 1799 771
rect 1903 209 1955 771
<< metal2 >>
rect 14 515 2284 771
rect 14 209 2284 465
<< labels >>
rlabel metal2 s 14 515 2284 771 6 DRAIN
port 1 nsew
rlabel metal1 s 381 843 1917 980 6 GATE
port 2 nsew
rlabel metal1 s 381 0 1917 137 6 GATE
port 2 nsew
rlabel metal2 s 14 209 2284 465 6 SOURCE
port 3 nsew
rlabel metal1 s 41 209 100 771 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 2198 209 2257 771 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 14 0 2284 980
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8649522
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8608492
string device primitive
<< end >>
