magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -36 679 4508 1471
<< pwell >>
rect 4336 25 4438 159
<< psubdiff >>
rect 4362 109 4412 133
rect 4362 75 4370 109
rect 4404 75 4412 109
rect 4362 51 4412 75
<< nsubdiff >>
rect 4362 1339 4412 1363
rect 4362 1305 4370 1339
rect 4404 1305 4412 1339
rect 4362 1281 4412 1305
<< psubdiffcont >>
rect 4370 75 4404 109
<< nsubdiffcont >>
rect 4370 1305 4404 1339
<< poly >>
rect 114 740 144 907
rect 48 724 144 740
rect 48 690 64 724
rect 98 690 144 724
rect 48 674 144 690
rect 114 507 144 674
<< polycont >>
rect 64 690 98 724
<< locali >>
rect 0 1397 4472 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 490 1130 524 1397
rect 706 1130 740 1397
rect 922 1130 956 1397
rect 1138 1130 1172 1397
rect 1354 1130 1388 1397
rect 1570 1130 1604 1397
rect 1786 1130 1820 1397
rect 2002 1130 2036 1397
rect 2218 1130 2252 1397
rect 2434 1130 2468 1397
rect 2650 1130 2684 1397
rect 2866 1130 2900 1397
rect 3082 1130 3116 1397
rect 3298 1130 3332 1397
rect 3514 1130 3548 1397
rect 3730 1130 3764 1397
rect 3946 1130 3980 1397
rect 4162 1130 4196 1397
rect 4370 1339 4404 1397
rect 4370 1289 4404 1305
rect 64 724 98 740
rect 64 674 98 690
rect 2216 724 2250 1096
rect 2216 690 2267 724
rect 2216 318 2250 690
rect 62 17 96 218
rect 274 17 308 218
rect 490 17 524 218
rect 706 17 740 218
rect 922 17 956 218
rect 1138 17 1172 218
rect 1354 17 1388 218
rect 1570 17 1604 218
rect 1786 17 1820 218
rect 2002 17 2036 218
rect 2218 17 2252 218
rect 2434 17 2468 218
rect 2650 17 2684 218
rect 2866 17 2900 218
rect 3082 17 3116 218
rect 3298 17 3332 218
rect 3514 17 3548 218
rect 3730 17 3764 218
rect 3946 17 3980 218
rect 4162 17 4196 218
rect 4370 109 4404 125
rect 4370 17 4404 75
rect 0 -17 4472 17
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_16  sky130_sram_1kbyte_1rw1r_32x256_8_contact_16_0
timestamp 1683767628
transform 1 0 48 0 1 674
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_28  sky130_sram_1kbyte_1rw1r_32x256_8_contact_28_0
timestamp 1683767628
transform 1 0 4362 0 1 1281
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_29  sky130_sram_1kbyte_1rw1r_32x256_8_contact_29_0
timestamp 1683767628
transform 1 0 4362 0 1 51
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m39_w2_000_sli_dli_da_p  sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m39_w2_000_sli_dli_da_p_0
timestamp 1683767628
transform 1 0 54 0 1 51
box -26 -26 4280 456
use sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m39_w2_000_sli_dli_da_p  sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m39_w2_000_sli_dli_da_p_0
timestamp 1683767628
transform 1 0 54 0 1 963
box -59 -56 4313 454
<< labels >>
rlabel locali s 81 707 81 707 4 A
rlabel locali s 2250 707 2250 707 4 Z
rlabel locali s 2236 0 2236 0 4 gnd
rlabel locali s 2236 1414 2236 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 4472 1414
string GDS_END 350156
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 345854
<< end >>
