magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 642 200 912 207
rect 454 191 912 200
rect 266 157 912 191
rect 1527 203 1711 207
rect 1527 157 1931 203
rect 1 71 1931 157
rect 1 64 640 71
rect 1 55 452 64
rect 1 21 353 55
rect 912 21 1931 71
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 247 47 277 131
rect 344 81 374 165
rect 532 90 562 174
rect 720 97 750 181
rect 804 97 834 181
rect 990 47 1020 131
rect 1074 47 1104 131
rect 1262 47 1292 131
rect 1450 47 1480 131
rect 1603 97 1633 181
rect 1823 47 1853 177
<< scpmoshvt >>
rect 79 413 109 497
rect 163 413 193 497
rect 351 363 381 447
rect 435 363 465 447
rect 623 413 653 497
rect 809 363 839 447
rect 893 363 923 447
rect 988 413 1018 497
rect 1072 413 1102 497
rect 1260 413 1290 497
rect 1448 413 1478 497
rect 1545 366 1575 450
rect 1823 297 1853 497
<< ndiff >>
rect 292 153 344 165
rect 292 131 300 153
rect 27 102 79 131
rect 27 68 35 102
rect 69 68 79 102
rect 27 47 79 68
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 47 247 131
rect 277 119 300 131
rect 334 119 344 153
rect 277 81 344 119
rect 374 127 426 165
rect 374 93 384 127
rect 418 93 426 127
rect 374 81 426 93
rect 480 136 532 174
rect 480 102 488 136
rect 522 102 532 136
rect 480 90 532 102
rect 562 145 614 174
rect 562 111 572 145
rect 606 111 614 145
rect 562 90 614 111
rect 668 143 720 181
rect 668 109 676 143
rect 710 109 720 143
rect 668 97 720 109
rect 750 169 804 181
rect 750 135 760 169
rect 794 135 804 169
rect 750 97 804 135
rect 834 169 886 181
rect 834 135 844 169
rect 878 135 886 169
rect 834 122 886 135
rect 1553 131 1603 181
rect 834 97 884 122
rect 940 105 990 131
rect 277 47 327 81
rect 938 93 990 105
rect 938 59 946 93
rect 980 59 990 93
rect 938 47 990 59
rect 1020 93 1074 131
rect 1020 59 1030 93
rect 1064 59 1074 93
rect 1020 47 1074 59
rect 1104 109 1156 131
rect 1104 75 1114 109
rect 1148 75 1156 109
rect 1104 47 1156 75
rect 1210 93 1262 131
rect 1210 59 1218 93
rect 1252 59 1262 93
rect 1210 47 1262 59
rect 1292 115 1344 131
rect 1292 81 1302 115
rect 1336 81 1344 115
rect 1292 47 1344 81
rect 1398 101 1450 131
rect 1398 67 1406 101
rect 1440 67 1450 101
rect 1398 47 1450 67
rect 1480 101 1603 131
rect 1480 67 1546 101
rect 1580 97 1603 101
rect 1633 169 1685 181
rect 1633 135 1643 169
rect 1677 135 1685 169
rect 1633 97 1685 135
rect 1580 67 1588 97
rect 1480 47 1588 67
rect 1771 93 1823 177
rect 1771 59 1779 93
rect 1813 59 1823 93
rect 1771 47 1823 59
rect 1853 101 1905 177
rect 1853 67 1863 101
rect 1897 67 1905 101
rect 1853 47 1905 67
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 413 79 443
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 413 163 451
rect 193 477 245 497
rect 193 443 203 477
rect 237 443 245 477
rect 571 477 623 497
rect 193 413 245 443
rect 299 409 351 447
rect 299 375 307 409
rect 341 375 351 409
rect 299 363 351 375
rect 381 425 435 447
rect 381 391 391 425
rect 425 391 435 425
rect 381 363 435 391
rect 465 421 515 447
rect 571 443 579 477
rect 613 443 623 477
rect 571 431 623 443
rect 465 409 517 421
rect 573 413 623 431
rect 653 485 705 497
rect 653 451 663 485
rect 697 451 705 485
rect 653 439 705 451
rect 938 447 988 497
rect 653 413 703 439
rect 759 421 809 447
rect 465 375 475 409
rect 509 375 517 409
rect 465 363 517 375
rect 757 409 809 421
rect 757 375 765 409
rect 799 375 809 409
rect 757 363 809 375
rect 839 425 893 447
rect 839 391 849 425
rect 883 391 893 425
rect 839 363 893 391
rect 923 413 988 447
rect 1018 485 1072 497
rect 1018 451 1028 485
rect 1062 451 1072 485
rect 1018 413 1072 451
rect 1102 477 1154 497
rect 1102 443 1112 477
rect 1146 443 1154 477
rect 1102 413 1154 443
rect 1208 485 1260 497
rect 1208 451 1216 485
rect 1250 451 1260 485
rect 1208 413 1260 451
rect 1290 477 1342 497
rect 1290 443 1300 477
rect 1334 443 1342 477
rect 1290 413 1342 443
rect 1396 477 1448 497
rect 1396 443 1404 477
rect 1438 443 1448 477
rect 1396 413 1448 443
rect 1478 485 1530 497
rect 1478 451 1488 485
rect 1522 451 1530 485
rect 1478 450 1530 451
rect 1771 485 1823 497
rect 1771 451 1779 485
rect 1813 451 1823 485
rect 1478 413 1545 450
rect 923 363 973 413
rect 1493 366 1545 413
rect 1575 425 1703 450
rect 1575 391 1585 425
rect 1619 391 1703 425
rect 1575 366 1703 391
rect 1771 297 1823 451
rect 1853 477 1905 497
rect 1853 443 1863 477
rect 1897 443 1905 477
rect 1853 297 1905 443
<< ndiffc >>
rect 35 68 69 102
rect 119 59 153 93
rect 300 119 334 153
rect 384 93 418 127
rect 488 102 522 136
rect 572 111 606 145
rect 676 109 710 143
rect 760 135 794 169
rect 844 135 878 169
rect 946 59 980 93
rect 1030 59 1064 93
rect 1114 75 1148 109
rect 1218 59 1252 93
rect 1302 81 1336 115
rect 1406 67 1440 101
rect 1546 67 1580 101
rect 1643 135 1677 169
rect 1779 59 1813 93
rect 1863 67 1897 101
<< pdiffc >>
rect 35 443 69 477
rect 119 451 153 485
rect 203 443 237 477
rect 307 375 341 409
rect 391 391 425 425
rect 579 443 613 477
rect 663 451 697 485
rect 475 375 509 409
rect 765 375 799 409
rect 849 391 883 425
rect 1028 451 1062 485
rect 1112 443 1146 477
rect 1216 451 1250 485
rect 1300 443 1334 477
rect 1404 443 1438 477
rect 1488 451 1522 485
rect 1779 451 1813 485
rect 1585 391 1619 425
rect 1863 443 1897 477
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 351 447 381 523
rect 435 447 465 523
rect 623 497 653 523
rect 79 265 109 413
rect 163 265 193 413
rect 809 447 839 523
rect 893 447 923 522
rect 988 497 1018 523
rect 1072 497 1102 523
rect 1260 497 1290 523
rect 1448 497 1478 523
rect 351 267 381 363
rect 435 348 465 363
rect 623 348 653 413
rect 1545 450 1575 523
rect 1823 497 1853 523
rect 809 348 839 363
rect 435 318 839 348
rect 532 273 645 318
rect 55 249 109 265
rect 55 215 65 249
rect 99 215 109 249
rect 55 199 109 215
rect 151 249 205 265
rect 151 215 161 249
rect 195 215 205 249
rect 151 199 205 215
rect 247 257 482 267
rect 247 237 432 257
rect 79 131 109 199
rect 163 131 193 199
rect 247 131 277 237
rect 416 223 432 237
rect 466 223 482 257
rect 416 213 482 223
rect 532 253 750 273
rect 893 265 923 363
rect 988 277 1018 413
rect 1072 277 1102 413
rect 532 219 666 253
rect 700 219 750 253
rect 532 199 750 219
rect 344 165 374 191
rect 532 174 562 199
rect 720 181 750 199
rect 804 253 923 265
rect 804 219 831 253
rect 865 235 923 253
rect 965 261 1030 277
rect 865 219 881 235
rect 804 209 881 219
rect 965 227 975 261
rect 1009 227 1030 261
rect 965 211 1030 227
rect 1072 261 1126 277
rect 1260 265 1290 413
rect 1448 265 1478 413
rect 1545 265 1575 366
rect 1823 265 1853 297
rect 1072 227 1082 261
rect 1116 227 1126 261
rect 1072 211 1126 227
rect 1201 249 1480 265
rect 1201 215 1211 249
rect 1245 215 1480 249
rect 1545 255 1704 265
rect 1545 235 1654 255
rect 804 181 834 209
rect 990 131 1020 211
rect 1074 131 1104 211
rect 1201 200 1480 215
rect 1201 199 1292 200
rect 1262 131 1292 199
rect 1450 131 1480 200
rect 1603 221 1654 235
rect 1688 221 1704 255
rect 1603 211 1704 221
rect 1779 249 1853 265
rect 1779 215 1791 249
rect 1825 215 1853 249
rect 1603 181 1633 211
rect 1779 199 1853 215
rect 344 51 374 81
rect 532 51 562 90
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 344 21 562 51
rect 720 21 750 97
rect 804 21 834 97
rect 1823 177 1853 199
rect 990 21 1020 47
rect 1074 21 1104 47
rect 1262 21 1292 47
rect 1450 21 1480 47
rect 1603 21 1633 97
rect 1823 21 1853 47
<< polycont >>
rect 65 215 99 249
rect 161 215 195 249
rect 432 223 466 257
rect 666 219 700 253
rect 831 219 865 253
rect 975 227 1009 261
rect 1082 227 1116 261
rect 1211 215 1245 249
rect 1654 221 1688 255
rect 1791 215 1825 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 35 477 69 493
rect 103 485 169 527
rect 103 451 119 485
rect 153 451 169 485
rect 203 477 509 493
rect 35 393 69 443
rect 237 459 509 477
rect 203 427 237 443
rect 307 409 341 425
rect 35 375 307 393
rect 35 359 341 375
rect 375 391 391 425
rect 425 391 441 425
rect 475 409 509 459
rect 375 325 409 391
rect 475 359 509 375
rect 543 477 613 493
rect 543 443 579 477
rect 647 485 713 527
rect 647 451 663 485
rect 697 451 713 485
rect 765 459 967 493
rect 543 325 613 443
rect 765 409 799 459
rect 30 249 99 323
rect 30 215 65 249
rect 30 199 99 215
rect 161 249 248 323
rect 195 215 248 249
rect 161 199 248 215
rect 282 291 409 325
rect 282 187 316 291
rect 452 279 613 325
rect 452 257 524 279
rect 416 223 432 257
rect 466 255 524 257
rect 466 223 490 255
rect 416 221 490 223
rect 35 127 237 161
rect 35 102 69 127
rect 35 52 69 68
rect 103 59 119 93
rect 153 59 169 93
rect 103 17 169 59
rect 203 85 237 127
rect 282 153 306 187
rect 282 119 300 153
rect 334 119 350 153
rect 384 127 418 152
rect 384 85 418 93
rect 452 136 524 221
rect 653 253 713 399
rect 765 357 799 375
rect 833 391 849 425
rect 883 391 899 425
rect 833 357 865 391
rect 933 417 967 459
rect 1012 485 1078 527
rect 1012 451 1028 485
rect 1062 451 1078 485
rect 1112 477 1146 493
rect 1196 485 1266 527
rect 1196 451 1216 485
rect 1250 451 1266 485
rect 1300 477 1337 493
rect 1112 417 1146 443
rect 1334 443 1337 477
rect 1300 427 1337 443
rect 933 383 1146 417
rect 833 323 899 357
rect 653 219 666 253
rect 700 219 713 253
rect 653 199 713 219
rect 747 289 899 323
rect 747 184 781 289
rect 960 261 1009 335
rect 815 219 831 253
rect 960 227 975 261
rect 865 219 881 221
rect 960 211 1009 227
rect 1050 261 1116 335
rect 1050 227 1082 261
rect 1050 211 1116 227
rect 1211 249 1269 335
rect 1245 215 1269 249
rect 1211 199 1269 215
rect 1303 255 1337 427
rect 1396 477 1438 493
rect 1396 443 1404 477
rect 1472 485 1729 493
rect 1472 451 1488 485
rect 1522 459 1729 485
rect 1522 451 1538 459
rect 1396 427 1438 443
rect 1303 221 1327 255
rect 747 169 810 184
rect 452 102 488 136
rect 522 102 524 136
rect 452 86 524 102
rect 560 145 618 161
rect 560 111 572 145
rect 606 111 618 145
rect 203 51 418 85
rect 560 17 618 111
rect 676 143 710 159
rect 744 135 760 169
rect 794 135 810 169
rect 744 119 810 135
rect 844 177 878 185
rect 844 169 1148 177
rect 878 143 1148 169
rect 844 119 878 135
rect 1099 109 1148 143
rect 1303 131 1337 221
rect 1396 187 1430 427
rect 1569 397 1585 425
rect 1478 391 1585 397
rect 1619 391 1635 425
rect 1478 357 1511 391
rect 1545 357 1635 391
rect 1478 351 1635 357
rect 1695 367 1729 459
rect 1763 485 1829 527
rect 1763 451 1779 485
rect 1813 451 1829 485
rect 1863 477 1915 493
rect 1897 443 1915 477
rect 1396 153 1410 187
rect 676 85 710 109
rect 1030 93 1064 109
rect 925 85 946 93
rect 676 59 946 85
rect 980 59 996 93
rect 676 51 996 59
rect 1099 75 1114 109
rect 1302 115 1337 131
rect 1478 117 1512 351
rect 1695 333 1825 367
rect 1638 221 1654 255
rect 1688 221 1695 255
rect 1791 249 1825 333
rect 1628 185 1676 187
rect 1628 169 1677 185
rect 1791 177 1825 215
rect 1628 153 1643 169
rect 1642 135 1643 153
rect 1642 119 1677 135
rect 1711 143 1825 177
rect 1099 59 1148 75
rect 1202 59 1218 93
rect 1252 59 1268 93
rect 1336 81 1337 115
rect 1302 65 1337 81
rect 1406 101 1512 117
rect 1440 83 1512 101
rect 1546 101 1580 117
rect 1030 17 1064 59
rect 1202 17 1268 59
rect 1406 51 1440 67
rect 1711 85 1745 143
rect 1580 67 1745 85
rect 1546 51 1745 67
rect 1779 93 1813 109
rect 1779 17 1813 59
rect 1863 101 1915 443
rect 1897 67 1915 101
rect 1863 51 1915 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 490 221 524 255
rect 306 153 340 187
rect 865 357 899 391
rect 858 253 892 255
rect 858 221 865 253
rect 865 221 892 253
rect 1327 221 1361 255
rect 1511 357 1545 391
rect 1410 153 1444 187
rect 1695 221 1729 255
rect 1594 153 1628 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 853 391 911 397
rect 853 357 865 391
rect 899 388 911 391
rect 1499 391 1557 397
rect 1499 388 1511 391
rect 899 360 1511 388
rect 899 357 911 360
rect 853 351 911 357
rect 1499 357 1511 360
rect 1545 357 1557 391
rect 1499 351 1557 357
rect 478 255 536 261
rect 478 221 490 255
rect 524 252 536 255
rect 846 255 904 261
rect 846 252 858 255
rect 524 224 858 252
rect 524 221 536 224
rect 478 215 536 221
rect 846 221 858 224
rect 892 221 904 255
rect 846 215 904 221
rect 1315 255 1373 261
rect 1315 221 1327 255
rect 1361 252 1373 255
rect 1683 255 1741 261
rect 1683 252 1695 255
rect 1361 224 1695 252
rect 1361 221 1373 224
rect 1315 215 1373 221
rect 1683 221 1695 224
rect 1729 221 1741 255
rect 1683 215 1741 221
rect 294 187 352 193
rect 294 153 306 187
rect 340 184 352 187
rect 1398 187 1456 193
rect 1398 184 1410 187
rect 340 156 1410 184
rect 340 153 352 156
rect 294 147 352 153
rect 1398 153 1410 156
rect 1444 184 1456 187
rect 1582 187 1640 193
rect 1582 184 1594 187
rect 1444 156 1594 184
rect 1444 153 1456 156
rect 1398 147 1456 153
rect 1582 153 1594 156
rect 1628 153 1640 187
rect 1582 147 1640 153
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
flabel locali s 674 289 708 323 0 FreeSans 200 0 0 0 S0
port 5 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A1
port 2 nsew signal input
flabel locali s 1870 221 1904 255 0 FreeSans 200 0 0 0 X
port 11 nsew signal output
flabel locali s 1870 289 1904 323 0 FreeSans 200 0 0 0 X
port 11 nsew signal output
flabel locali s 1870 357 1904 391 0 FreeSans 200 0 0 0 X
port 11 nsew signal output
flabel locali s 1235 221 1269 255 0 FreeSans 200 0 0 0 S1
port 6 nsew signal input
flabel locali s 1057 221 1091 255 0 FreeSans 200 0 0 0 A2
port 3 nsew signal input
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 A1
port 2 nsew signal input
flabel locali s 214 289 248 323 0 FreeSans 200 0 0 0 A0
port 1 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 A0
port 1 nsew signal input
flabel locali s 1870 153 1904 187 0 FreeSans 200 0 0 0 X
port 11 nsew signal output
flabel locali s 960 221 994 255 0 FreeSans 200 0 0 0 A3
port 4 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 8 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 9 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 7 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 10 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 mux4_1
rlabel metal1 s 0 -48 1932 48 1 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1932 592 1 VPWR
port 10 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1932 544
string GDS_END 1770002
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1754526
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 48.300 0.000 
<< end >>
