magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< pwell >>
rect -26 -26 176 98
<< scnmos >>
rect 60 0 90 72
<< ndiff >>
rect 0 53 60 72
rect 0 19 8 53
rect 42 19 60 53
rect 0 0 60 19
rect 90 53 150 72
rect 90 19 108 53
rect 142 19 150 53
rect 90 0 150 19
<< ndiffc >>
rect 8 19 42 53
rect 108 19 142 53
<< poly >>
rect 60 72 90 98
rect 60 -26 90 0
<< locali >>
rect 8 53 42 69
rect 8 3 42 19
rect 108 53 142 69
rect 108 3 142 19
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_11  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_11_0
timestamp 1683767628
transform 1 0 100 0 1 3
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_11  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_11_1
timestamp 1683767628
transform 1 0 0 0 1 3
box 0 0 1 1
<< labels >>
rlabel locali s 25 36 25 36 4 S
rlabel locali s 125 36 125 36 4 D
rlabel poly s 75 36 75 36 4 G
<< properties >>
string FIXED_BBOX -25 -26 175 98
string GDS_END 1950
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 1154
<< end >>
