magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< locali >>
rect 169 1140 177 1174
rect 211 1140 249 1174
rect 283 1140 321 1174
rect 355 1140 393 1174
rect 427 1140 465 1174
rect 499 1140 507 1174
rect 169 20 177 54
rect 211 20 249 54
rect 283 20 321 54
rect 355 20 393 54
rect 427 20 465 54
rect 499 20 507 54
<< viali >>
rect 177 1140 211 1174
rect 249 1140 283 1174
rect 321 1140 355 1174
rect 393 1140 427 1174
rect 465 1140 499 1174
rect 177 20 211 54
rect 249 20 283 54
rect 321 20 355 54
rect 393 20 427 54
rect 465 20 499 54
<< obsli1 >>
rect 38 1010 72 1048
rect 38 938 72 976
rect 38 866 72 904
rect 38 794 72 832
rect 38 722 72 760
rect 38 650 72 688
rect 38 578 72 616
rect 38 506 72 544
rect 38 434 72 472
rect 38 362 72 400
rect 38 290 72 328
rect 38 218 72 256
rect 38 112 72 184
rect 149 88 183 1106
rect 235 88 269 1106
rect 321 88 355 1106
rect 407 88 441 1106
rect 493 88 527 1106
rect 604 1010 638 1048
rect 604 938 638 976
rect 604 866 638 904
rect 604 794 638 832
rect 604 722 638 760
rect 604 650 638 688
rect 604 578 638 616
rect 604 506 638 544
rect 604 434 638 472
rect 604 362 638 400
rect 604 290 638 328
rect 604 218 638 256
rect 604 112 638 184
<< obsli1c >>
rect 38 1048 72 1082
rect 38 976 72 1010
rect 38 904 72 938
rect 38 832 72 866
rect 38 760 72 794
rect 38 688 72 722
rect 38 616 72 650
rect 38 544 72 578
rect 38 472 72 506
rect 38 400 72 434
rect 38 328 72 362
rect 38 256 72 290
rect 38 184 72 218
rect 604 1048 638 1082
rect 604 976 638 1010
rect 604 904 638 938
rect 604 832 638 866
rect 604 760 638 794
rect 604 688 638 722
rect 604 616 638 650
rect 604 544 638 578
rect 604 472 638 506
rect 604 400 638 434
rect 604 328 638 362
rect 604 256 638 290
rect 604 184 638 218
<< metal1 >>
rect 165 1174 511 1194
rect 165 1140 177 1174
rect 211 1140 249 1174
rect 283 1140 321 1174
rect 355 1140 393 1174
rect 427 1140 465 1174
rect 499 1140 511 1174
rect 165 1128 511 1140
rect 26 1082 84 1094
rect 26 1048 38 1082
rect 72 1048 84 1082
rect 26 1010 84 1048
rect 26 976 38 1010
rect 72 976 84 1010
rect 26 938 84 976
rect 26 904 38 938
rect 72 904 84 938
rect 26 866 84 904
rect 26 832 38 866
rect 72 832 84 866
rect 26 794 84 832
rect 26 760 38 794
rect 72 760 84 794
rect 26 722 84 760
rect 26 688 38 722
rect 72 688 84 722
rect 26 650 84 688
rect 26 616 38 650
rect 72 616 84 650
rect 26 578 84 616
rect 26 544 38 578
rect 72 544 84 578
rect 26 506 84 544
rect 26 472 38 506
rect 72 472 84 506
rect 26 434 84 472
rect 26 400 38 434
rect 72 400 84 434
rect 26 362 84 400
rect 26 328 38 362
rect 72 328 84 362
rect 26 290 84 328
rect 26 256 38 290
rect 72 256 84 290
rect 26 218 84 256
rect 26 184 38 218
rect 72 184 84 218
rect 26 100 84 184
rect 592 1082 650 1094
rect 592 1048 604 1082
rect 638 1048 650 1082
rect 592 1010 650 1048
rect 592 976 604 1010
rect 638 976 650 1010
rect 592 938 650 976
rect 592 904 604 938
rect 638 904 650 938
rect 592 866 650 904
rect 592 832 604 866
rect 638 832 650 866
rect 592 794 650 832
rect 592 760 604 794
rect 638 760 650 794
rect 592 722 650 760
rect 592 688 604 722
rect 638 688 650 722
rect 592 650 650 688
rect 592 616 604 650
rect 638 616 650 650
rect 592 578 650 616
rect 592 544 604 578
rect 638 544 650 578
rect 592 506 650 544
rect 592 472 604 506
rect 638 472 650 506
rect 592 434 650 472
rect 592 400 604 434
rect 638 400 650 434
rect 592 362 650 400
rect 592 328 604 362
rect 638 328 650 362
rect 592 290 650 328
rect 592 256 604 290
rect 638 256 650 290
rect 592 218 650 256
rect 592 184 604 218
rect 638 184 650 218
rect 592 100 650 184
rect 165 54 511 66
rect 165 20 177 54
rect 211 20 249 54
rect 283 20 321 54
rect 355 20 393 54
rect 427 20 465 54
rect 499 20 511 54
rect 165 0 511 20
<< obsm1 >>
rect 140 100 192 1094
rect 226 100 278 1094
rect 312 100 364 1094
rect 398 100 450 1094
rect 484 100 536 1094
<< metal2 >>
rect 0 622 676 1094
rect 0 100 676 572
<< labels >>
rlabel metal2 s 0 622 676 1094 6 DRAIN
port 1 nsew
rlabel viali s 465 1140 499 1174 6 GATE
port 2 nsew
rlabel viali s 465 20 499 54 6 GATE
port 2 nsew
rlabel viali s 393 1140 427 1174 6 GATE
port 2 nsew
rlabel viali s 393 20 427 54 6 GATE
port 2 nsew
rlabel viali s 321 1140 355 1174 6 GATE
port 2 nsew
rlabel viali s 321 20 355 54 6 GATE
port 2 nsew
rlabel viali s 249 1140 283 1174 6 GATE
port 2 nsew
rlabel viali s 249 20 283 54 6 GATE
port 2 nsew
rlabel viali s 177 1140 211 1174 6 GATE
port 2 nsew
rlabel viali s 177 20 211 54 6 GATE
port 2 nsew
rlabel locali s 169 1140 507 1174 6 GATE
port 2 nsew
rlabel locali s 169 20 507 54 6 GATE
port 2 nsew
rlabel metal1 s 165 1128 511 1194 6 GATE
port 2 nsew
rlabel metal1 s 165 0 511 66 6 GATE
port 2 nsew
rlabel metal2 s 0 100 676 572 6 SOURCE
port 3 nsew
rlabel metal1 s 26 100 84 1094 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 592 100 650 1094 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 676 1194
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6138690
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 6116728
<< end >>
