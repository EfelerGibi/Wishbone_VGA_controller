magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1 201 1637 203
rect 1 23 1951 201
rect 1 21 479 23
rect 956 21 1140 23
rect 1552 21 1951 23
rect 47 -17 81 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 468 93 498 177
rect 662 49 692 177
rect 772 49 802 177
rect 1034 47 1064 177
rect 1220 49 1250 177
rect 1372 49 1402 133
rect 1531 49 1561 177
rect 1651 47 1681 167
rect 1751 47 1781 175
rect 1843 47 1873 175
<< scpmoshvt >>
rect 99 297 129 497
rect 183 297 213 497
rect 267 297 297 497
rect 351 297 381 497
rect 450 297 480 425
rect 654 325 684 493
rect 760 325 790 493
rect 1001 297 1031 497
rect 1220 297 1250 465
rect 1372 297 1402 425
rect 1547 329 1577 457
rect 1650 329 1680 497
rect 1751 297 1781 497
rect 1843 297 1873 497
<< ndiff >>
rect 27 93 79 177
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 129 163 177
rect 109 95 119 129
rect 153 95 163 129
rect 109 47 163 95
rect 193 93 247 177
rect 193 59 203 93
rect 237 59 247 93
rect 193 47 247 59
rect 277 129 331 177
rect 277 95 287 129
rect 321 95 331 129
rect 277 47 331 95
rect 361 93 468 177
rect 498 169 554 177
rect 498 135 508 169
rect 542 135 554 169
rect 498 93 554 135
rect 608 165 662 177
rect 608 131 618 165
rect 652 131 662 165
rect 361 89 453 93
rect 361 55 371 89
rect 405 55 453 89
rect 361 47 453 55
rect 608 49 662 131
rect 692 91 772 177
rect 692 57 702 91
rect 736 57 772 91
rect 692 49 772 57
rect 802 169 901 177
rect 802 135 854 169
rect 888 135 901 169
rect 802 49 901 135
rect 982 161 1034 177
rect 982 127 990 161
rect 1024 127 1034 161
rect 982 93 1034 127
rect 982 59 990 93
rect 1024 59 1034 93
rect 982 47 1034 59
rect 1064 161 1116 177
rect 1064 127 1074 161
rect 1108 127 1116 161
rect 1064 121 1116 127
rect 1064 47 1114 121
rect 1170 105 1220 177
rect 1168 97 1220 105
rect 1168 63 1176 97
rect 1210 63 1220 97
rect 1168 49 1220 63
rect 1250 133 1351 177
rect 1427 169 1531 177
rect 1427 135 1473 169
rect 1507 135 1531 169
rect 1427 133 1531 135
rect 1250 126 1372 133
rect 1250 92 1260 126
rect 1294 92 1372 126
rect 1250 49 1372 92
rect 1402 49 1531 133
rect 1561 167 1611 177
rect 1701 167 1751 175
rect 1561 93 1651 167
rect 1561 59 1573 93
rect 1607 59 1651 93
rect 1561 49 1651 59
rect 1578 47 1651 49
rect 1681 142 1751 167
rect 1681 108 1707 142
rect 1741 108 1751 142
rect 1681 47 1751 108
rect 1781 97 1843 175
rect 1781 63 1799 97
rect 1833 63 1843 97
rect 1781 47 1843 63
rect 1873 101 1925 175
rect 1873 67 1883 101
rect 1917 67 1925 101
rect 1873 47 1925 67
<< pdiff >>
rect 47 477 99 497
rect 47 443 55 477
rect 89 443 99 477
rect 47 297 99 443
rect 129 477 183 497
rect 129 443 139 477
rect 173 443 183 477
rect 129 409 183 443
rect 129 375 139 409
rect 173 375 183 409
rect 129 341 183 375
rect 129 307 139 341
rect 173 307 183 341
rect 129 297 183 307
rect 213 477 267 497
rect 213 443 223 477
rect 257 443 267 477
rect 213 297 267 443
rect 297 477 351 497
rect 297 443 307 477
rect 341 443 351 477
rect 297 409 351 443
rect 297 375 307 409
rect 341 375 351 409
rect 297 341 351 375
rect 297 307 307 341
rect 341 307 351 341
rect 297 297 351 307
rect 381 477 433 497
rect 381 443 391 477
rect 425 443 433 477
rect 381 425 433 443
rect 381 297 450 425
rect 480 341 544 425
rect 480 307 498 341
rect 532 307 544 341
rect 602 413 654 493
rect 602 379 610 413
rect 644 379 654 413
rect 602 325 654 379
rect 684 481 760 493
rect 684 447 703 481
rect 737 447 760 481
rect 684 325 760 447
rect 790 481 895 493
rect 790 447 850 481
rect 884 447 895 481
rect 790 325 895 447
rect 949 481 1001 497
rect 949 447 957 481
rect 991 447 1001 481
rect 480 297 544 307
rect 949 297 1001 447
rect 1031 349 1081 497
rect 1135 405 1220 465
rect 1135 371 1143 405
rect 1177 371 1220 405
rect 1135 365 1220 371
rect 1031 343 1083 349
rect 1031 309 1041 343
rect 1075 309 1083 343
rect 1031 297 1083 309
rect 1137 297 1220 365
rect 1250 425 1350 465
rect 1592 489 1650 497
rect 1592 457 1604 489
rect 1462 425 1547 457
rect 1250 409 1372 425
rect 1250 375 1301 409
rect 1335 375 1372 409
rect 1250 341 1372 375
rect 1250 307 1301 341
rect 1335 307 1372 341
rect 1250 297 1372 307
rect 1402 421 1547 425
rect 1402 387 1503 421
rect 1537 387 1547 421
rect 1402 329 1547 387
rect 1577 455 1604 457
rect 1638 455 1650 489
rect 1577 329 1650 455
rect 1680 341 1751 497
rect 1680 329 1707 341
rect 1402 297 1497 329
rect 1695 307 1707 329
rect 1741 307 1751 341
rect 1695 297 1751 307
rect 1781 489 1843 497
rect 1781 455 1799 489
rect 1833 455 1843 489
rect 1781 297 1843 455
rect 1873 477 1925 497
rect 1873 443 1883 477
rect 1917 443 1925 477
rect 1873 409 1925 443
rect 1873 375 1883 409
rect 1917 375 1925 409
rect 1873 297 1925 375
<< ndiffc >>
rect 35 59 69 93
rect 119 95 153 129
rect 203 59 237 93
rect 287 95 321 129
rect 508 135 542 169
rect 618 131 652 165
rect 371 55 405 89
rect 702 57 736 91
rect 854 135 888 169
rect 990 127 1024 161
rect 990 59 1024 93
rect 1074 127 1108 161
rect 1176 63 1210 97
rect 1473 135 1507 169
rect 1260 92 1294 126
rect 1573 59 1607 93
rect 1707 108 1741 142
rect 1799 63 1833 97
rect 1883 67 1917 101
<< pdiffc >>
rect 55 443 89 477
rect 139 443 173 477
rect 139 375 173 409
rect 139 307 173 341
rect 223 443 257 477
rect 307 443 341 477
rect 307 375 341 409
rect 307 307 341 341
rect 391 443 425 477
rect 498 307 532 341
rect 610 379 644 413
rect 703 447 737 481
rect 850 447 884 481
rect 957 447 991 481
rect 1143 371 1177 405
rect 1041 309 1075 343
rect 1301 375 1335 409
rect 1301 307 1335 341
rect 1503 387 1537 421
rect 1604 455 1638 489
rect 1707 307 1741 341
rect 1799 455 1833 489
rect 1883 443 1917 477
rect 1883 375 1917 409
<< poly >>
rect 99 497 129 523
rect 183 497 213 523
rect 267 497 297 523
rect 351 497 381 523
rect 654 493 684 519
rect 760 493 790 519
rect 1001 497 1031 523
rect 450 425 480 483
rect 99 265 129 297
rect 183 265 213 297
rect 267 265 297 297
rect 351 265 381 297
rect 450 265 480 297
rect 654 271 684 325
rect 654 265 693 271
rect 760 265 790 325
rect 1220 493 1577 523
rect 1650 497 1680 523
rect 1751 497 1781 523
rect 1843 497 1873 523
rect 1220 465 1250 493
rect 1547 457 1577 493
rect 1372 425 1402 451
rect 80 249 408 265
rect 80 215 364 249
rect 398 215 408 249
rect 80 207 408 215
rect 79 199 408 207
rect 450 249 693 265
rect 450 215 581 249
rect 615 215 649 249
rect 683 215 693 249
rect 450 199 693 215
rect 748 249 802 265
rect 748 215 758 249
rect 792 215 802 249
rect 1001 247 1031 297
rect 1220 247 1250 297
rect 1372 265 1402 297
rect 1547 265 1577 329
rect 1001 217 1250 247
rect 748 199 802 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 331 177 361 199
rect 468 177 498 199
rect 662 197 693 199
rect 662 177 692 197
rect 772 177 802 199
rect 1034 177 1064 217
rect 1220 177 1250 217
rect 1292 249 1402 265
rect 1292 215 1302 249
rect 1336 215 1402 249
rect 1292 199 1402 215
rect 468 67 498 93
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 662 21 692 49
rect 772 21 802 49
rect 1372 133 1402 199
rect 1531 249 1585 265
rect 1650 256 1680 329
rect 1751 265 1781 297
rect 1843 265 1873 297
rect 1650 255 1681 256
rect 1531 215 1541 249
rect 1575 215 1585 249
rect 1531 199 1585 215
rect 1627 239 1681 255
rect 1627 205 1637 239
rect 1671 205 1681 239
rect 1531 177 1561 199
rect 1627 189 1681 205
rect 1723 249 1781 265
rect 1723 215 1733 249
rect 1767 215 1781 249
rect 1723 199 1781 215
rect 1823 249 1877 265
rect 1823 215 1833 249
rect 1867 215 1877 249
rect 1823 199 1877 215
rect 1651 167 1681 189
rect 1751 175 1781 199
rect 1843 175 1873 199
rect 1034 21 1064 47
rect 1220 21 1250 49
rect 1372 23 1402 49
rect 1531 21 1561 49
rect 1651 21 1681 47
rect 1751 21 1781 47
rect 1843 21 1873 47
<< polycont >>
rect 364 215 398 249
rect 581 215 615 249
rect 649 215 683 249
rect 758 215 792 249
rect 1302 215 1336 249
rect 1541 215 1575 249
rect 1637 205 1671 239
rect 1733 215 1767 249
rect 1833 215 1867 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 55 477 89 527
rect 55 427 89 443
rect 139 477 173 493
rect 207 477 273 527
rect 207 443 223 477
rect 257 443 273 477
rect 307 477 341 493
rect 375 477 441 527
rect 941 481 1007 527
rect 1783 489 1849 527
rect 375 443 391 477
rect 425 443 441 477
rect 475 447 703 481
rect 737 447 783 481
rect 826 447 850 481
rect 884 447 907 481
rect 941 447 957 481
rect 991 447 1007 481
rect 1074 455 1604 489
rect 1638 455 1693 489
rect 1783 455 1799 489
rect 1833 455 1849 489
rect 1883 477 1935 493
rect 139 409 173 443
rect 307 409 341 443
rect 475 409 509 447
rect 873 413 907 447
rect 1074 413 1108 455
rect 173 375 307 409
rect 139 341 341 375
rect 173 307 307 341
rect 139 291 341 307
rect 375 375 509 409
rect 578 379 610 413
rect 644 379 839 413
rect 873 379 1108 413
rect 1143 405 1177 421
rect 139 288 284 291
rect 221 185 284 288
rect 375 265 409 375
rect 474 307 498 341
rect 532 307 771 341
rect 364 249 409 265
rect 398 215 409 249
rect 364 193 409 215
rect 119 166 307 185
rect 375 173 409 193
rect 119 132 321 166
rect 375 139 473 173
rect 119 129 153 132
rect 35 93 69 109
rect 119 70 153 95
rect 287 129 321 132
rect 35 17 69 59
rect 187 59 203 93
rect 237 59 253 93
rect 287 70 321 95
rect 371 89 405 105
rect 187 17 253 59
rect 371 17 405 55
rect 439 85 473 139
rect 508 169 542 307
rect 737 265 771 307
rect 805 339 839 379
rect 805 323 911 339
rect 805 305 877 323
rect 854 289 877 305
rect 854 275 911 289
rect 576 249 703 265
rect 576 215 581 249
rect 615 215 649 249
rect 683 215 703 249
rect 576 199 703 215
rect 737 249 811 265
rect 737 215 758 249
rect 792 215 811 249
rect 737 199 811 215
rect 854 169 888 275
rect 945 241 979 379
rect 1025 309 1041 343
rect 1075 309 1108 343
rect 1025 289 1108 309
rect 508 119 542 135
rect 598 131 618 165
rect 652 131 820 165
rect 682 85 702 91
rect 439 57 702 85
rect 736 57 752 91
rect 439 51 752 57
rect 786 85 820 131
rect 854 119 888 135
rect 922 210 979 241
rect 922 209 978 210
rect 922 208 976 209
rect 922 207 973 208
rect 922 85 956 207
rect 1060 187 1108 289
rect 786 51 956 85
rect 990 161 1024 177
rect 990 93 1024 127
rect 1060 153 1061 187
rect 1095 161 1108 187
rect 1060 127 1074 153
rect 1060 83 1108 127
rect 1143 119 1177 371
rect 1215 178 1249 455
rect 1917 443 1935 477
rect 1883 421 1935 443
rect 1283 375 1301 409
rect 1335 375 1366 409
rect 1283 341 1366 375
rect 1283 307 1301 341
rect 1335 323 1366 341
rect 1473 387 1503 421
rect 1537 409 1935 421
rect 1537 387 1883 409
rect 1335 307 1337 323
rect 1283 289 1337 307
rect 1371 289 1439 323
rect 1286 249 1371 254
rect 1286 215 1302 249
rect 1336 215 1371 249
rect 1286 199 1371 215
rect 1328 187 1371 199
rect 1215 165 1255 178
rect 1215 144 1294 165
rect 1221 131 1294 144
rect 1260 126 1294 131
rect 1328 153 1337 187
rect 1328 126 1371 153
rect 1143 85 1153 119
rect 990 17 1024 59
rect 1143 63 1176 85
rect 1210 63 1226 97
rect 1260 64 1294 92
rect 1405 85 1439 289
rect 1473 169 1507 387
rect 1838 375 1883 387
rect 1917 375 1935 409
rect 1541 289 1657 323
rect 1691 307 1707 341
rect 1741 307 1855 341
rect 1691 299 1855 307
rect 1541 249 1575 289
rect 1821 265 1855 299
rect 1541 199 1575 215
rect 1609 239 1671 255
rect 1609 205 1637 239
rect 1705 249 1787 265
rect 1705 215 1733 249
rect 1767 215 1787 249
rect 1821 249 1867 265
rect 1821 215 1833 249
rect 1609 189 1671 205
rect 1821 199 1867 215
rect 1609 187 1650 189
rect 1609 153 1613 187
rect 1647 153 1650 187
rect 1821 181 1855 199
rect 1609 146 1650 153
rect 1707 150 1855 181
rect 1699 147 1855 150
rect 1473 119 1507 135
rect 1699 142 1757 147
rect 1699 119 1707 142
rect 1541 85 1573 93
rect 1143 53 1226 63
rect 1405 59 1573 85
rect 1607 59 1634 93
rect 1699 85 1705 119
rect 1741 108 1757 142
rect 1901 117 1935 375
rect 1739 85 1757 108
rect 1699 59 1757 85
rect 1799 97 1833 113
rect 1405 51 1634 59
rect 1799 17 1833 63
rect 1883 101 1935 117
rect 1917 67 1935 101
rect 1883 51 1935 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 877 289 911 323
rect 1061 161 1095 187
rect 1061 153 1074 161
rect 1074 153 1095 161
rect 1337 289 1371 323
rect 1337 153 1371 187
rect 1153 97 1187 119
rect 1153 85 1176 97
rect 1176 85 1187 97
rect 1613 153 1647 187
rect 1705 108 1707 119
rect 1707 108 1739 119
rect 1705 85 1739 108
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 865 323 923 329
rect 865 289 877 323
rect 911 320 923 323
rect 1325 323 1383 329
rect 1325 320 1337 323
rect 911 292 1337 320
rect 911 289 923 292
rect 865 283 923 289
rect 1325 289 1337 292
rect 1371 289 1383 323
rect 1325 283 1383 289
rect 1049 187 1107 193
rect 1049 153 1061 187
rect 1095 184 1107 187
rect 1325 187 1383 193
rect 1325 184 1337 187
rect 1095 156 1337 184
rect 1095 153 1107 156
rect 1049 147 1107 153
rect 1325 153 1337 156
rect 1371 184 1383 187
rect 1601 187 1659 193
rect 1601 184 1613 187
rect 1371 156 1613 184
rect 1371 153 1383 156
rect 1325 147 1383 153
rect 1601 153 1613 156
rect 1647 153 1659 187
rect 1601 147 1659 153
rect 1141 119 1199 125
rect 1141 85 1153 119
rect 1187 116 1199 119
rect 1693 119 1751 125
rect 1693 116 1705 119
rect 1187 88 1705 116
rect 1187 85 1199 88
rect 1141 79 1199 85
rect 1693 85 1705 88
rect 1739 85 1751 119
rect 1693 79 1751 85
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
flabel locali s 233 357 267 391 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 601 221 635 255 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1613 289 1647 323 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1705 221 1739 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel pwell s 47 -17 81 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 47 527 81 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 1799 17 1833 113 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel locali s 1783 455 1849 527 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 hkscl5hdv1_xor3_1
flabel comment s 0 544 0 544 3 FreeSans 200 0 0 0 HHNEC
rlabel locali s 990 17 1024 177 1 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 371 17 405 105 1 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 187 17 253 93 1 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 35 17 69 109 1 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 0 -17 2024 17 1 VGND
port 4 nsew ground bidirectional abutment
rlabel locali s 941 447 1007 527 1 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 375 443 441 527 1 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 207 443 273 527 1 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 55 427 89 527 1 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 0 527 2024 561 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2024 544
string GDS_END 698948
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 685650
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 10.120 0.000 
<< end >>
