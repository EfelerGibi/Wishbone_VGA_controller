magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< obsm2 >>
rect -6231 21500 -1085 23500
tri -1915 21330 -1745 21500 ne
rect -1745 21330 -1085 21500
tri -1085 21330 1085 23500 sw
tri -1745 18500 1085 21330 ne
tri 1085 20500 1915 21330 sw
rect 1085 18500 6008 20500
rect -6231 15500 -1085 17500
tri -1915 15330 -1745 15500 ne
rect -1745 15330 -1085 15500
tri -1085 15330 1085 17500 sw
tri -1745 12500 1085 15330 ne
tri 1085 14500 1915 15330 sw
rect 1085 12500 6008 14500
rect 9908 -1000 27500 1000
tri -915 -17500 1085 -15500 se
rect 1085 -17500 6008 -15500
tri -1915 -18500 -915 -17500 se
rect -915 -18500 915 -17500
tri 915 -18500 1915 -17500 nw
rect -6231 -20500 -1085 -18500
tri -1085 -20500 915 -18500 nw
tri -915 -23500 1085 -21500 se
rect 1085 -23500 6008 -21500
tri -1915 -24500 -915 -23500 se
rect -915 -24500 915 -23500
tri 915 -24500 1915 -23500 nw
rect -6231 -26500 -1085 -24500
tri -1085 -26500 915 -24500 nw
<< obsm3 >>
tri -13806 23672 -10978 26500 se
rect -10978 24500 10978 26500
tri -10978 23672 -10150 24500 nw
tri 10150 23672 10978 24500 ne
tri 10978 23672 13806 26500 sw
tri -16634 20844 -13806 23672 se
rect -13806 22290 -12360 23672
tri -12360 22290 -10978 23672 nw
tri -10946 22290 -9736 23500 se
rect -9736 23253 -2202 23500
tri -2202 23253 -1955 23500 sw
rect -9736 22290 -1955 23253
rect -13806 22104 -12546 22290
tri -12546 22104 -12360 22290 nw
tri -11132 22104 -10946 22290 se
rect -10946 22104 -1955 22290
tri -13806 20844 -12546 22104 nw
tri -12392 20844 -11132 22104 se
rect -11132 21747 -1955 22104
tri -668 21747 1085 23500 se
rect 1085 22290 9736 23500
tri 9736 22290 10946 23500 sw
tri 10978 22290 12360 23672 ne
rect 12360 23500 13806 23672
tri 13806 23500 13978 23672 sw
rect 12360 22290 13978 23500
rect 1085 21747 10946 22290
rect -11132 21500 -2202 21747
tri -2202 21500 -1955 21747 nw
rect -11132 20844 -9736 21500
tri -19462 18016 -16634 20844 se
rect -16634 19895 -14755 20844
tri -14755 19895 -13806 20844 nw
tri -13341 19895 -12392 20844 se
rect -12392 20672 -9736 20844
tri -9736 20672 -8908 21500 nw
rect -12392 19895 -10513 20672
tri -10513 19895 -9736 20672 nw
tri -1915 20500 -668 21747 se
rect -668 21500 10946 21747
rect -668 20500 915 21500
tri 915 20500 1915 21500 nw
tri -9098 19895 -8493 20500 se
rect -8493 20151 566 20500
tri 566 20151 915 20500 nw
tri 1732 20253 1979 20500 se
rect 1979 20253 8493 20500
rect 1732 20151 8493 20253
tri 8493 20151 8842 20500 sw
tri 8908 20151 10257 21500 ne
rect 10257 21048 10946 21500
tri 10946 21048 12188 22290 sw
tri 12360 21048 13602 22290 ne
rect 13602 21048 13978 22290
tri 13978 21048 16430 23500 sw
rect 10257 20151 12188 21048
rect -8493 19895 -738 20151
rect -16634 19371 -15279 19895
tri -15279 19371 -14755 19895 nw
tri -13865 19371 -13341 19895 se
rect -13341 19371 -11305 19895
tri -16634 18016 -15279 19371 nw
tri -15220 18016 -13865 19371 se
rect -13865 19103 -11305 19371
tri -11305 19103 -10513 19895 nw
tri -9890 19103 -9098 19895 se
rect -9098 19103 -738 19895
rect -13865 18016 -12564 19103
tri -22290 15188 -19462 18016 se
rect -19462 16629 -18021 18016
tri -18021 16629 -16634 18016 nw
tri -16607 16629 -15220 18016 se
rect -15220 17844 -12564 18016
tri -12564 17844 -11305 19103 nw
tri -11149 17844 -9890 19103 se
rect -9890 18847 -738 19103
tri -738 18847 566 20151 nw
rect -9890 18500 -1085 18847
tri -1085 18500 -738 18847 nw
rect 1732 18747 8842 20151
tri 8842 18747 10246 20151 sw
tri 10257 18747 11661 20151 ne
rect 11661 19634 12188 20151
tri 12188 19634 13602 21048 sw
tri 13602 19634 15016 21048 ne
rect 15016 19634 16430 21048
tri 16430 19634 17844 21048 sw
rect 11661 18747 13602 19634
tri 1732 18500 1979 18747 ne
rect 1979 18500 10246 18747
tri 10246 18500 10493 18747 sw
tri 11661 18500 11908 18747 ne
rect 11908 18500 13602 18747
rect -9890 17844 -8493 18500
rect -15220 16629 -13978 17844
rect -19462 16430 -18220 16629
tri -18220 16430 -18021 16629 nw
tri -16806 16430 -16607 16629 se
rect -16607 16430 -13978 16629
tri -13978 16430 -12564 17844 nw
tri -12563 16430 -11149 17844 se
rect -11149 17672 -8493 17844
tri -8493 17672 -7665 18500 nw
rect -11149 16430 -9906 17672
tri -19462 15188 -18220 16430 nw
tri -23849 13629 -22290 15188 se
rect -22290 15016 -19634 15188
tri -19634 15016 -19462 15188 nw
tri -18220 15016 -16806 16430 se
rect -16806 16373 -14035 16430
tri -14035 16373 -13978 16430 nw
tri -12620 16373 -12563 16430 se
rect -12563 16373 -9906 16430
rect -16806 15016 -15392 16373
tri -15392 15016 -14035 16373 nw
tri -13977 15016 -12620 16373 se
rect -12620 16259 -9906 16373
tri -9906 16259 -8493 17672 nw
tri -8492 16259 -7251 17500 se
rect -7251 17253 -2202 17500
tri -2202 17253 -1955 17500 sw
rect -7251 16259 -1955 17253
rect -12620 16105 -10060 16259
tri -10060 16105 -9906 16259 nw
tri -8646 16105 -8492 16259 se
rect -8492 16105 -1955 16259
rect -12620 15016 -11321 16105
rect -22290 13629 -21021 15016
tri -21021 13629 -19634 15016 nw
tri -19607 13629 -18220 15016 se
rect -18220 13629 -16806 15016
tri -26500 10978 -23849 13629 se
rect -23849 12360 -22290 13629
tri -22290 12360 -21021 13629 nw
tri -20876 12360 -19607 13629 se
rect -19607 13602 -16806 13629
tri -16806 13602 -15392 15016 nw
tri -15391 13602 -13977 15016 se
rect -13977 14844 -11321 15016
tri -11321 14844 -10060 16105 nw
tri -9907 14844 -8646 16105 se
rect -8646 15747 -1955 16105
tri -668 15747 1085 17500 se
rect 1085 17149 7251 17500
tri 7251 17149 7602 17500 sw
tri 7665 17149 9016 18500 ne
rect 9016 17149 10493 18500
tri 10493 17149 11844 18500 sw
tri 11908 17149 13259 18500 ne
rect 13259 18220 13602 18500
tri 13602 18220 15016 19634 sw
tri 15016 18220 16430 19634 ne
rect 16430 18220 17844 19634
rect 13259 17149 15016 18220
rect 1085 15747 7602 17149
rect -8646 15500 -2202 15747
tri -2202 15500 -1955 15747 nw
rect -8646 14844 -7251 15500
rect -13977 13602 -12734 14844
rect -19607 12360 -18220 13602
rect -23849 10978 -23672 12360
tri -23672 10978 -22290 12360 nw
tri -22258 10978 -20876 12360 se
rect -20876 12188 -18220 12360
tri -18220 12188 -16806 13602 nw
tri -16805 12188 -15391 13602 se
rect -15391 13431 -12734 13602
tri -12734 13431 -11321 14844 nw
tri -11320 13431 -9907 14844 se
rect -9907 14672 -7251 14844
tri -7251 14672 -6423 15500 nw
rect -9907 13431 -8665 14672
rect -15391 13373 -12792 13431
tri -12792 13373 -12734 13431 nw
tri -11378 13373 -11320 13431 se
rect -11320 13373 -8665 13431
rect -15391 12188 -14149 13373
rect -20876 10978 -19430 12188
tri -19430 10978 -18220 12188 nw
tri -18015 10978 -16805 12188 se
rect -16805 12016 -14149 12188
tri -14149 12016 -12792 13373 nw
tri -12735 12016 -11378 13373 se
rect -11378 13258 -8665 13373
tri -8665 13258 -7251 14672 nw
tri -1915 14500 -668 15747 se
rect -668 15735 7602 15747
tri 7602 15735 9016 17149 sw
tri 9016 15735 10430 17149 ne
rect 10430 15735 11844 17149
tri 11844 15735 13258 17149 sw
tri 13259 15735 14673 17149 ne
rect 14673 16806 15016 17149
tri 15016 16806 16430 18220 sw
tri 16430 16806 17844 18220 ne
tri 17844 16806 20672 19634 sw
rect 14673 15735 16430 16806
rect -668 15500 9016 15735
rect -668 14500 915 15500
tri 915 14500 1915 15500 nw
tri -7250 13258 -6008 14500 se
rect -6008 14149 564 14500
tri 564 14149 915 14500 nw
tri 1732 14253 1979 14500 se
rect 1979 14253 6008 14500
rect 1732 14149 6008 14253
tri 6008 14149 6359 14500 sw
tri 6423 14149 7774 15500 ne
rect 7774 14321 9016 15500
tri 9016 14321 10430 15735 sw
tri 10430 14321 11844 15735 ne
rect 11844 14321 13258 15735
tri 13258 14321 14672 15735 sw
tri 14673 14321 16087 15735 ne
rect 16087 15392 16430 15735
tri 16430 15392 17844 16806 sw
tri 17844 15392 19258 16806 ne
rect 19258 15392 20672 16806
rect 16087 14321 17844 15392
rect 7774 14149 10430 14321
rect -6008 13258 -736 14149
rect -11378 13105 -8818 13258
tri -8818 13105 -8665 13258 nw
tri -7403 13105 -7250 13258 se
rect -7250 13105 -736 13258
rect -11378 12016 -10079 13105
rect -16805 10978 -15562 12016
rect -26500 -10978 -24500 10978
tri -24500 10150 -23672 10978 nw
tri -23500 9736 -22258 10978 se
rect -22258 9736 -20672 10978
tri -20672 9736 -19430 10978 nw
tri -19257 9736 -18015 10978 se
rect -18015 10603 -15562 10978
tri -15562 10603 -14149 12016 nw
tri -14148 10603 -12735 12016 se
rect -12735 11844 -10079 12016
tri -10079 11844 -8818 13105 nw
tri -8664 11844 -7403 13105 se
rect -7403 12849 -736 13105
tri -736 12849 564 14149 nw
rect -7403 12500 -1085 12849
tri -1085 12500 -736 12849 nw
rect 1732 12747 6359 14149
tri 6359 12747 7761 14149 sw
tri 7774 12747 9176 14149 ne
rect 9176 12907 10430 14149
tri 10430 12907 11844 14321 sw
tri 11844 12907 13258 14321 ne
rect 13258 12907 14672 14321
tri 14672 12907 16086 14321 sw
tri 16087 12907 17501 14321 ne
rect 17501 13978 17844 14321
tri 17844 13978 19258 15392 sw
tri 19258 13978 20672 15392 ne
tri 20672 13978 23500 16806 sw
rect 17501 12907 19258 13978
rect 9176 12747 11844 12907
tri 1732 12500 1979 12747 ne
rect 1979 12500 7761 12747
tri 7761 12500 8008 12747 sw
tri 9176 12500 9423 12747 ne
rect 9423 12500 11844 12747
rect -7403 11844 -6016 12500
rect -12735 10603 -11493 11844
rect -18015 10430 -15735 10603
tri -15735 10430 -15562 10603 nw
tri -14321 10430 -14148 10603 se
rect -14148 10430 -11493 10603
tri -11493 10430 -10079 11844 nw
tri -10078 10430 -8664 11844 se
rect -8664 11664 -6016 11844
tri -6016 11664 -5180 12500 nw
rect -8664 10430 -7421 11664
rect -18015 9736 -16977 10430
rect -23500 -9736 -21500 9736
tri -21500 8908 -20672 9736 nw
tri -20500 8493 -19257 9736 se
rect -19257 9188 -16977 9736
tri -16977 9188 -15735 10430 nw
tri -15563 9188 -14321 10430 se
rect -14321 9188 -12907 10430
rect -19257 8493 -17672 9188
tri -17672 8493 -16977 9188 nw
tri -16258 8493 -15563 9188 se
rect -15563 9016 -12907 9188
tri -12907 9016 -11493 10430 nw
tri -11492 9016 -10078 10430 se
rect -10078 10259 -7421 10430
tri -7421 10259 -6016 11664 nw
rect -10078 9016 -8836 10259
rect -15563 8908 -13015 9016
tri -13015 8908 -12907 9016 nw
tri -11600 8908 -11492 9016 se
rect -11492 8908 -8836 9016
rect -15563 8493 -14258 8908
rect -20500 -8493 -18500 8493
tri -18500 7665 -17672 8493 nw
tri -17500 7251 -16258 8493 se
rect -16258 7665 -14258 8493
tri -14258 7665 -13015 8908 nw
tri -12843 7665 -11600 8908 se
rect -11600 8844 -8836 8908
tri -8836 8844 -7421 10259 nw
tri 5180 10079 7601 12500 ne
rect 7601 11664 8008 12500
tri 8008 11664 8844 12500 sw
tri 9423 11664 10259 12500 ne
rect 10259 11664 11844 12500
rect 7601 10251 8844 11664
tri 8844 10251 10257 11664 sw
tri 10259 10251 11672 11664 ne
rect 11672 11493 11844 11664
tri 11844 11493 13258 12907 sw
tri 13258 11493 14672 12907 ne
rect 14672 11493 16086 12907
tri 16086 11493 17500 12907 sw
tri 17501 11493 18915 12907 ne
rect 18915 12564 19258 12907
tri 19258 12564 20672 13978 sw
tri 20672 12564 22086 13978 ne
rect 22086 12564 23500 13978
rect 18915 11493 20672 12564
rect 11672 10251 13258 11493
rect 7601 10079 10257 10251
tri 7601 8844 8836 10079 ne
rect 8836 8844 10257 10079
rect -11600 7665 -11257 8844
rect -16258 7251 -15500 7665
rect -17500 -7251 -15500 7251
tri -15500 6423 -14258 7665 nw
tri -14085 6423 -12843 7665 se
rect -12843 6423 -11257 7665
tri -11257 6423 -8836 8844 nw
tri 8836 7431 10249 8844 ne
rect 10249 8836 10257 8844
tri 10257 8836 11672 10251 sw
tri 11672 10079 11844 10251 ne
rect 11844 10079 13258 10251
tri 13258 10079 14672 11493 sw
tri 14672 10079 16086 11493 ne
rect 16086 10079 17500 11493
tri 17500 10079 18914 11493 sw
tri 18915 10079 20329 11493 ne
rect 20329 11150 20672 11493
tri 20672 11150 22086 12564 sw
tri 22086 11150 23500 12564 ne
tri 23500 11150 26328 13978 sw
rect 20329 10079 22086 11150
tri 11844 8836 13087 10079 ne
rect 13087 8836 14672 10079
rect 10249 7431 11672 8836
tri 10249 6423 11257 7431 ne
rect 11257 7423 11672 7431
tri 11672 7423 13085 8836 sw
tri 13087 7665 14258 8836 ne
rect 14258 8665 14672 8836
tri 14672 8665 16086 10079 sw
tri 16086 8665 17500 10079 ne
rect 17500 8665 18914 10079
tri 18914 8665 20328 10079 sw
tri 20329 8908 21500 10079 ne
rect 21500 9736 22086 10079
tri 22086 9736 23500 11150 sw
tri 23500 10150 24500 11150 ne
rect 24500 10978 26328 11150
tri 26328 10978 26500 11150 sw
rect 14258 7665 16086 8665
tri 14258 7423 14500 7665 ne
rect 14500 7423 16086 7665
rect 11257 6423 13085 7423
tri -14500 6008 -14085 6423 se
rect -14085 6008 -12500 6423
rect -14500 1000 -12500 6008
tri -12500 5180 -11257 6423 nw
tri 11257 5180 12500 6423 ne
rect 12500 6008 13085 6423
tri 13085 6008 14500 7423 sw
tri 14500 6423 15500 7423 ne
rect 15500 7251 16086 7423
tri 16086 7251 17500 8665 sw
tri 17500 7665 18500 8665 ne
rect 18500 8493 20328 8665
tri 20328 8493 20500 8665 sw
rect -14500 -1000 11500 1000
rect -14500 -6008 -12500 -1000
tri -14500 -6423 -14085 -6008 ne
rect -14085 -6423 -12500 -6008
tri -17500 -7665 -17086 -7251 ne
rect -17086 -7665 -15500 -7251
tri -15500 -7665 -14258 -6423 sw
tri -14085 -7665 -12843 -6423 ne
rect -12843 -7665 -12500 -6423
tri -12500 -7665 -10015 -5180 sw
tri 10257 -7423 12500 -5180 se
rect 12500 -6008 14500 6008
rect 12500 -7251 13257 -6008
tri 13257 -7251 14500 -6008 nw
tri 14672 -7251 15500 -6423 se
rect 15500 -7251 17500 7251
rect 12500 -7423 12843 -7251
tri -20500 -8908 -20085 -8493 ne
rect -20085 -8908 -18500 -8493
tri -18500 -8908 -17257 -7665 sw
tri -17086 -8908 -15843 -7665 ne
rect -15843 -8665 -14258 -7665
tri -14258 -8665 -13258 -7665 sw
tri -12843 -8665 -11843 -7665 ne
rect -11843 -8665 -10015 -7665
rect -15843 -8908 -13258 -8665
tri -26500 -12360 -25118 -10978 ne
rect -25118 -11150 -24500 -10978
tri -24500 -11150 -23500 -10150 sw
tri -23500 -11150 -22086 -9736 ne
rect -22086 -10150 -21500 -9736
tri -21500 -10150 -20258 -8908 sw
tri -20085 -10150 -18843 -8908 ne
rect -18843 -9908 -17257 -8908
tri -17257 -9908 -16257 -8908 sw
tri -15843 -9908 -14843 -8908 ne
rect -14843 -9908 -13258 -8908
rect -18843 -10150 -16257 -9908
rect -22086 -11150 -20258 -10150
tri -20258 -11150 -19258 -10150 sw
tri -18843 -11150 -17843 -10150 ne
rect -17843 -11150 -16257 -10150
rect -25118 -12360 -23500 -11150
tri -25118 -13806 -23672 -12360 ne
rect -23672 -12564 -23500 -12360
tri -23500 -12564 -22086 -11150 sw
tri -22086 -12564 -20672 -11150 ne
rect -20672 -12564 -19258 -11150
tri -19258 -12564 -17844 -11150 sw
tri -17843 -11321 -17672 -11150 ne
rect -17672 -11321 -16257 -11150
tri -16257 -11321 -14844 -9908 sw
tri -14843 -10079 -14672 -9908 ne
rect -14672 -10079 -13258 -9908
tri -13258 -10079 -11844 -8665 sw
tri -11843 -10079 -10429 -8665 ne
rect -10429 -10079 -10015 -8665
tri -17672 -12564 -16429 -11321 ne
rect -16429 -11493 -14844 -11321
tri -14844 -11493 -14672 -11321 sw
tri -14672 -11493 -13258 -10079 ne
rect -13258 -11493 -11844 -10079
tri -11844 -11493 -10430 -10079 sw
tri -10429 -10251 -10257 -10079 ne
rect -10257 -10251 -10015 -10079
tri -10015 -10251 -7429 -7665 sw
tri 7601 -10079 10257 -7423 se
rect 10257 -7665 12843 -7423
tri 12843 -7665 13257 -7251 nw
rect 10257 -8493 12015 -7665
tri 12015 -8493 12843 -7665 nw
tri 13430 -8493 14672 -7251 se
rect 14672 -8493 16086 -7251
rect 10257 -9736 10772 -8493
tri 10772 -9736 12015 -8493 nw
tri 12187 -9736 13430 -8493 se
rect 13430 -8665 16086 -8493
tri 16086 -8665 17500 -7251 nw
tri 17500 -8665 18500 -7665 se
rect 18500 -8493 20500 8493
rect 18500 -8665 19257 -8493
rect 13430 -9736 14672 -8665
rect 10257 -10079 10358 -9736
tri -10257 -11493 -9015 -10251 ne
rect -9015 -11493 -7429 -10251
rect -16429 -12564 -14672 -11493
rect -23672 -13806 -22086 -12564
tri -23672 -15188 -22290 -13806 ne
rect -22290 -13978 -22086 -13806
tri -22086 -13978 -20672 -12564 sw
tri -20672 -13978 -19258 -12564 ne
rect -19258 -13978 -17844 -12564
tri -17844 -13978 -16430 -12564 sw
tri -16429 -13978 -15015 -12564 ne
rect -15015 -12907 -14672 -12564
tri -14672 -12907 -13258 -11493 sw
tri -13258 -12907 -11844 -11493 ne
rect -11844 -12907 -10430 -11493
tri -10430 -12907 -9016 -11493 sw
tri -9015 -12907 -7601 -11493 ne
rect -7601 -11664 -7429 -11493
tri -7429 -11664 -6016 -10251 sw
rect -7601 -12500 -6016 -11664
tri -6016 -12500 -5180 -11664 sw
tri 5180 -12500 7601 -10079 se
rect 7601 -10150 10358 -10079
tri 10358 -10150 10772 -9736 nw
tri 11773 -10150 12187 -9736 se
rect 12187 -10079 14672 -9736
tri 14672 -10079 16086 -8665 nw
tri 16086 -10079 17500 -8665 se
rect 17500 -9736 19257 -8665
tri 19257 -9736 20500 -8493 nw
tri 20672 -9736 21500 -8908 se
rect 21500 -9736 23500 9736
rect 24500 5000 26500 10978
rect 24500 3000 27500 5000
rect 17500 -10079 18015 -9736
rect 12187 -10150 14492 -10079
rect 7601 -11321 9187 -10150
tri 9187 -11321 10358 -10150 nw
tri 10602 -11321 11773 -10150 se
rect 11773 -10259 14492 -10150
tri 14492 -10259 14672 -10079 nw
tri 15906 -10259 16086 -10079 se
rect 16086 -10259 18015 -10079
rect 11773 -11321 13430 -10259
tri 13430 -11321 14492 -10259 nw
tri 14844 -11321 15906 -10259 se
rect 15906 -10978 18015 -10259
tri 18015 -10978 19257 -9736 nw
tri 19430 -10978 20672 -9736 se
rect 20672 -10978 22258 -9736
tri 22258 -10978 23500 -9736 nw
rect 24500 -5000 27500 -3000
tri 23672 -10978 24500 -10150 se
rect 24500 -10978 26500 -5000
rect 15906 -11321 16633 -10978
rect 7601 -12500 8008 -11321
tri 8008 -12500 9187 -11321 nw
tri 9423 -12500 10602 -11321 se
rect 10602 -12500 12187 -11321
rect -7601 -12907 6702 -12500
rect -15015 -13978 -13258 -12907
rect -22290 -15188 -20672 -13978
tri -22290 -16634 -20844 -15188 ne
rect -20844 -15392 -20672 -15188
tri -20672 -15392 -19258 -13978 sw
tri -19258 -15392 -17844 -13978 ne
rect -17844 -15392 -16430 -13978
tri -16430 -15392 -15016 -13978 sw
tri -15015 -15392 -13601 -13978 ne
rect -13601 -14321 -13258 -13978
tri -13258 -14321 -11844 -12907 sw
tri -11844 -14321 -10430 -12907 ne
rect -10430 -14321 -9016 -12907
tri -9016 -14321 -7602 -12907 sw
tri -7601 -14149 -6359 -12907 ne
rect -6359 -13806 6702 -12907
tri 6702 -13806 8008 -12500 nw
tri 8117 -13806 9423 -12500 se
rect 9423 -12564 12187 -12500
tri 12187 -12564 13430 -11321 nw
tri 13601 -12564 14844 -11321 se
rect 14844 -12360 16633 -11321
tri 16633 -12360 18015 -10978 nw
tri 18048 -12360 19430 -10978 se
rect 19430 -12360 20876 -10978
tri 20876 -12360 22258 -10978 nw
tri 22290 -12360 23672 -10978 se
rect 23672 -12360 23876 -10978
rect 14844 -12564 15735 -12360
rect 9423 -13087 11664 -12564
tri 11664 -13087 12187 -12564 nw
tri 13078 -13087 13601 -12564 se
rect 13601 -13087 15735 -12564
rect 9423 -13806 10251 -13087
rect -6359 -14149 6008 -13806
rect -13601 -15392 -11844 -14321
rect -20844 -16634 -19258 -15392
tri -20844 -18016 -19462 -16634 ne
rect -19462 -16806 -19258 -16634
tri -19258 -16806 -17844 -15392 sw
tri -17844 -16806 -16430 -15392 ne
rect -16430 -16806 -15016 -15392
tri -15016 -16806 -13602 -15392 sw
tri -13601 -16806 -12187 -15392 ne
rect -12187 -15735 -11844 -15392
tri -11844 -15735 -10430 -14321 sw
tri -10430 -15735 -9016 -14321 ne
rect -9016 -15500 -7602 -14321
tri -7602 -15500 -6423 -14321 sw
tri -6359 -14500 -6008 -14149 ne
rect -6008 -14500 6008 -14149
tri 6008 -14500 6702 -13806 nw
tri 7423 -14500 8117 -13806 se
rect 8117 -14500 10251 -13806
tri 10251 -14500 11664 -13087 nw
tri 11665 -14500 13078 -13087 se
rect 13078 -13258 15735 -13087
tri 15735 -13258 16633 -12360 nw
tri 17150 -13258 18048 -12360 se
rect 18048 -13258 19805 -12360
rect 13078 -14500 14321 -13258
tri 6423 -15500 7423 -14500 se
rect 7423 -15500 9004 -14500
rect -9016 -15735 -1085 -15500
rect -12187 -16806 -10430 -15735
rect -19462 -18016 -17844 -16806
tri -19462 -19628 -17850 -18016 ne
rect -17850 -18220 -17844 -18016
tri -17844 -18220 -16430 -16806 sw
tri -16430 -18220 -15016 -16806 ne
rect -15016 -18220 -13602 -16806
tri -13602 -18220 -12188 -16806 sw
tri -12187 -18220 -10773 -16806 ne
rect -10773 -17149 -10430 -16806
tri -10430 -17149 -9016 -15735 sw
tri -9016 -16977 -7774 -15735 ne
rect -7774 -16977 -1085 -15735
tri -7774 -17149 -7602 -16977 ne
rect -7602 -17149 -1085 -16977
rect -10773 -18220 -9016 -17149
rect -17850 -19628 -16430 -18220
tri -17850 -20844 -16634 -19628 ne
rect -16634 -19634 -16430 -19628
tri -16430 -19634 -15016 -18220 sw
tri -15016 -19634 -13602 -18220 ne
rect -13602 -19634 -12188 -18220
tri -12188 -19634 -10774 -18220 sw
tri -10773 -19634 -9359 -18220 ne
rect -9359 -18500 -9016 -18220
tri -9016 -18500 -7665 -17149 sw
tri -7602 -17500 -7251 -17149 ne
rect -7251 -17500 -1085 -17149
tri -1915 -18220 -1195 -17500 ne
rect -1195 -18220 -1085 -17500
tri -1085 -18220 1635 -15500 sw
tri 1732 -15747 1979 -15500 se
rect 1979 -15747 9004 -15500
tri 9004 -15747 10251 -14500 nw
tri 10418 -15747 11665 -14500 se
rect 11665 -14672 14321 -14500
tri 14321 -14672 15735 -13258 nw
tri 15736 -14672 17150 -13258 se
rect 17150 -13431 19805 -13258
tri 19805 -13431 20876 -12360 nw
tri 21219 -13431 22290 -12360 se
rect 22290 -13431 23876 -12360
rect 17150 -14672 18392 -13431
rect 11665 -15747 12907 -14672
rect 1732 -17149 7602 -15747
tri 7602 -17149 9004 -15747 nw
tri 9016 -17149 10418 -15747 se
rect 10418 -16086 12907 -15747
tri 12907 -16086 14321 -14672 nw
tri 14322 -16086 15736 -14672 se
rect 15736 -14844 18392 -14672
tri 18392 -14844 19805 -13431 nw
tri 19806 -14844 21219 -13431 se
rect 21219 -13602 23876 -13431
tri 23876 -13602 26500 -10978 nw
rect 21219 -14844 22462 -13602
rect 15736 -15016 18220 -14844
tri 18220 -15016 18392 -14844 nw
rect 15736 -16086 16977 -15016
rect 10418 -17149 11493 -16086
rect 1732 -17253 7498 -17149
tri 7498 -17253 7602 -17149 nw
tri 8912 -17253 9016 -17149 se
rect 9016 -17253 11493 -17149
tri 1732 -17500 1979 -17253 ne
rect 1979 -17500 7251 -17253
tri 7251 -17500 7498 -17253 nw
rect -9359 -18747 -2202 -18500
tri -2202 -18747 -1955 -18500 sw
rect -9359 -19634 -1955 -18747
rect -16634 -20844 -15016 -19634
tri -16634 -22372 -15106 -20844 ne
rect -15106 -21048 -15016 -20844
tri -15016 -21048 -13602 -19634 sw
tri -13602 -21048 -12188 -19634 ne
rect -12188 -21048 -10774 -19634
tri -10774 -21048 -9360 -19634 sw
tri -9359 -20500 -8493 -19634 ne
rect -8493 -20253 -1955 -19634
rect -8493 -20500 -2202 -20253
tri -2202 -20500 -1955 -20253 nw
tri -1195 -20500 1085 -18220 ne
rect 1085 -18500 1635 -18220
tri 1635 -18500 1915 -18220 sw
tri 7665 -18500 8912 -17253 se
rect 8912 -17500 11493 -17253
tri 11493 -17500 12907 -16086 nw
tri 12908 -17500 14322 -16086 se
rect 14322 -16259 16977 -16086
tri 16977 -16259 18220 -15016 nw
tri 19462 -15188 19806 -14844 se
rect 19806 -15016 22462 -14844
tri 22462 -15016 23876 -13602 nw
rect 19806 -15188 21048 -15016
tri 18391 -16259 19462 -15188 se
rect 19462 -16259 21048 -15188
rect 14322 -17500 15564 -16259
rect 8912 -18500 10493 -17500
tri 10493 -18500 11493 -17500 nw
tri 11908 -18500 12908 -17500 se
rect 12908 -17672 15564 -17500
tri 15564 -17672 16977 -16259 nw
tri 16978 -17672 18391 -16259 se
rect 18391 -16430 21048 -16259
tri 21048 -16430 22462 -15016 nw
rect 18391 -17672 19634 -16430
rect 12908 -17844 15392 -17672
tri 15392 -17844 15564 -17672 nw
rect 12908 -18500 14149 -17844
rect 1085 -19087 9906 -18500
tri 9906 -19087 10493 -18500 nw
tri 11321 -19087 11908 -18500 se
rect 11908 -19087 14149 -18500
tri 14149 -19087 15392 -17844 nw
tri 16634 -18016 16978 -17672 se
rect 16978 -17844 19634 -17672
tri 19634 -17844 21048 -16430 nw
rect 16978 -18016 18220 -17844
tri 15563 -19087 16634 -18016 se
rect 16634 -19087 18220 -18016
rect 1085 -20500 8493 -19087
tri 8493 -20500 9906 -19087 nw
tri 9908 -20500 11321 -19087 se
rect 11321 -20500 12736 -19087
tri 12736 -20500 14149 -19087 nw
tri 14150 -20500 15563 -19087 se
rect 15563 -19258 18220 -19087
tri 18220 -19258 19634 -17844 nw
rect 15563 -20500 16806 -19258
rect -15106 -22372 -13602 -21048
tri -15106 -23672 -13806 -22372 ne
rect -13806 -22462 -13602 -22372
tri -13602 -22462 -12188 -21048 sw
tri -12188 -22462 -10774 -21048 ne
rect -10774 -21500 -9360 -21048
tri -9360 -21500 -8908 -21048 sw
tri 8908 -21500 9908 -20500 se
rect 9908 -21500 11489 -20500
rect -10774 -22462 -1085 -21500
rect -13806 -23672 -12188 -22462
tri -12188 -23672 -10978 -22462 sw
tri -10774 -23500 -9736 -22462 ne
rect -9736 -23500 -1085 -22462
tri -1915 -23672 -1743 -23500 ne
rect -1743 -23672 -1085 -23500
tri -1085 -23672 1087 -21500 sw
tri 1732 -21747 1979 -21500 se
rect 1979 -21747 11489 -21500
tri 11489 -21747 12736 -20500 nw
tri 12903 -21747 14150 -20500 se
rect 14150 -20672 16806 -20500
tri 16806 -20672 18220 -19258 nw
rect 14150 -21747 15392 -20672
rect 1732 -22462 10774 -21747
tri 10774 -22462 11489 -21747 nw
tri 12188 -22462 12903 -21747 se
rect 12903 -22086 15392 -21747
tri 15392 -22086 16806 -20672 nw
rect 12903 -22462 13978 -22086
rect 1732 -23253 9983 -22462
tri 9983 -23253 10774 -22462 nw
tri 11397 -23253 12188 -22462 se
rect 12188 -23253 13978 -22462
tri 1732 -23500 1979 -23253 ne
rect 1979 -23500 9736 -23253
tri 9736 -23500 9983 -23253 nw
tri -13806 -26500 -10978 -23672 ne
tri -10978 -24500 -10150 -23672 sw
rect -10978 -24747 -2202 -24500
tri -2202 -24747 -1955 -24500 sw
rect -10978 -26253 -1955 -24747
rect -10978 -26500 -2202 -26253
tri -2202 -26500 -1955 -26253 nw
tri -1743 -26500 1085 -23672 ne
rect 1085 -24500 1087 -23672
tri 1087 -24500 1915 -23672 sw
tri 10150 -24500 11397 -23253 se
rect 11397 -23500 13978 -23253
tri 13978 -23500 15392 -22086 nw
rect 11397 -24500 12978 -23500
tri 12978 -24500 13978 -23500 nw
rect 1085 -26500 10978 -24500
tri 10978 -26500 12978 -24500 nw
<< properties >>
string FIXED_BBOX -26500 -26500 27500 26500
string LEFclass BLOCK
string LEFview TRUE
string gencell sky130_fd_pr__rf_test_coil2
string library sky130
string parameter m=1
string GDS_END 10411040
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10392572
<< end >>
