magic
tech sky130A
timestamp 1683767628
<< properties >>
string GDS_END 40006440
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 40005672
<< end >>
