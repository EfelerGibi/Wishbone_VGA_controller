magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -66 377 160 1251
rect 560 403 1054 863
rect 1454 493 2178 1251
rect 1960 377 2178 493
<< pwell >>
rect -26 1585 2138 1671
rect 668 1195 1394 1585
rect 1850 1345 2108 1585
rect 1174 317 1900 433
rect 600 43 1900 317
rect -26 -43 2138 43
<< mvnmos >>
rect 747 1221 847 1521
rect 903 1221 1003 1521
rect 1059 1221 1159 1521
rect 1215 1221 1315 1521
rect 1929 1371 2029 1521
rect 679 141 779 291
rect 835 141 935 291
rect 1253 107 1353 407
rect 1409 107 1509 407
rect 1565 107 1665 407
rect 1721 107 1821 407
<< mvpmos >>
rect 1593 885 1793 969
rect 1929 885 2029 1185
rect 679 469 779 619
rect 835 469 935 619
rect 1593 563 1793 647
<< mvndiff >>
rect 694 1509 747 1521
rect 694 1475 702 1509
rect 736 1475 747 1509
rect 694 1429 747 1475
rect 694 1395 702 1429
rect 736 1395 747 1429
rect 694 1347 747 1395
rect 694 1313 702 1347
rect 736 1313 747 1347
rect 694 1267 747 1313
rect 694 1233 702 1267
rect 736 1233 747 1267
rect 694 1221 747 1233
rect 847 1509 903 1521
rect 847 1475 858 1509
rect 892 1475 903 1509
rect 847 1429 903 1475
rect 847 1395 858 1429
rect 892 1395 903 1429
rect 847 1347 903 1395
rect 847 1313 858 1347
rect 892 1313 903 1347
rect 847 1267 903 1313
rect 847 1233 858 1267
rect 892 1233 903 1267
rect 847 1221 903 1233
rect 1003 1509 1059 1521
rect 1003 1475 1014 1509
rect 1048 1475 1059 1509
rect 1003 1429 1059 1475
rect 1003 1395 1014 1429
rect 1048 1395 1059 1429
rect 1003 1347 1059 1395
rect 1003 1313 1014 1347
rect 1048 1313 1059 1347
rect 1003 1267 1059 1313
rect 1003 1233 1014 1267
rect 1048 1233 1059 1267
rect 1003 1221 1059 1233
rect 1159 1509 1215 1521
rect 1159 1475 1170 1509
rect 1204 1475 1215 1509
rect 1159 1429 1215 1475
rect 1159 1395 1170 1429
rect 1204 1395 1215 1429
rect 1159 1347 1215 1395
rect 1159 1313 1170 1347
rect 1204 1313 1215 1347
rect 1159 1267 1215 1313
rect 1159 1233 1170 1267
rect 1204 1233 1215 1267
rect 1159 1221 1215 1233
rect 1315 1509 1368 1521
rect 1315 1475 1326 1509
rect 1360 1475 1368 1509
rect 1315 1429 1368 1475
rect 1315 1395 1326 1429
rect 1360 1395 1368 1429
rect 1315 1347 1368 1395
rect 1876 1509 1929 1521
rect 1876 1475 1884 1509
rect 1918 1475 1929 1509
rect 1876 1417 1929 1475
rect 1876 1383 1884 1417
rect 1918 1383 1929 1417
rect 1876 1371 1929 1383
rect 2029 1509 2082 1521
rect 2029 1475 2040 1509
rect 2074 1475 2082 1509
rect 2029 1417 2082 1475
rect 2029 1383 2040 1417
rect 2074 1383 2082 1417
rect 2029 1371 2082 1383
rect 1315 1313 1326 1347
rect 1360 1313 1368 1347
rect 1315 1267 1368 1313
rect 1315 1233 1326 1267
rect 1360 1233 1368 1267
rect 1315 1221 1368 1233
rect 1200 395 1253 407
rect 1200 361 1208 395
rect 1242 361 1253 395
rect 1200 315 1253 361
rect 626 279 679 291
rect 626 245 634 279
rect 668 245 679 279
rect 626 187 679 245
rect 626 153 634 187
rect 668 153 679 187
rect 626 141 679 153
rect 779 279 835 291
rect 779 245 790 279
rect 824 245 835 279
rect 779 187 835 245
rect 779 153 790 187
rect 824 153 835 187
rect 779 141 835 153
rect 935 279 988 291
rect 935 245 946 279
rect 980 245 988 279
rect 935 187 988 245
rect 935 153 946 187
rect 980 153 988 187
rect 935 141 988 153
rect 1200 281 1208 315
rect 1242 281 1253 315
rect 1200 233 1253 281
rect 1200 199 1208 233
rect 1242 199 1253 233
rect 1200 153 1253 199
rect 1200 119 1208 153
rect 1242 119 1253 153
rect 1200 107 1253 119
rect 1353 395 1409 407
rect 1353 361 1364 395
rect 1398 361 1409 395
rect 1353 315 1409 361
rect 1353 281 1364 315
rect 1398 281 1409 315
rect 1353 233 1409 281
rect 1353 199 1364 233
rect 1398 199 1409 233
rect 1353 153 1409 199
rect 1353 119 1364 153
rect 1398 119 1409 153
rect 1353 107 1409 119
rect 1509 395 1565 407
rect 1509 361 1520 395
rect 1554 361 1565 395
rect 1509 315 1565 361
rect 1509 281 1520 315
rect 1554 281 1565 315
rect 1509 233 1565 281
rect 1509 199 1520 233
rect 1554 199 1565 233
rect 1509 153 1565 199
rect 1509 119 1520 153
rect 1554 119 1565 153
rect 1509 107 1565 119
rect 1665 395 1721 407
rect 1665 361 1676 395
rect 1710 361 1721 395
rect 1665 315 1721 361
rect 1665 281 1676 315
rect 1710 281 1721 315
rect 1665 233 1721 281
rect 1665 199 1676 233
rect 1710 199 1721 233
rect 1665 153 1721 199
rect 1665 119 1676 153
rect 1710 119 1721 153
rect 1665 107 1721 119
rect 1821 395 1874 407
rect 1821 361 1832 395
rect 1866 361 1874 395
rect 1821 315 1874 361
rect 1821 281 1832 315
rect 1866 281 1874 315
rect 1821 233 1874 281
rect 1821 199 1832 233
rect 1866 199 1874 233
rect 1821 153 1874 199
rect 1821 119 1832 153
rect 1866 119 1874 153
rect 1821 107 1874 119
<< mvpdiff >>
rect 1520 999 1578 1011
rect 1520 965 1536 999
rect 1570 969 1578 999
rect 1876 1173 1929 1185
rect 1876 1139 1884 1173
rect 1918 1139 1929 1173
rect 1876 1093 1929 1139
rect 1876 1059 1884 1093
rect 1918 1059 1929 1093
rect 1876 1011 1929 1059
rect 1876 977 1884 1011
rect 1918 977 1929 1011
rect 1876 969 1929 977
rect 1570 965 1593 969
rect 1520 931 1593 965
rect 1520 897 1548 931
rect 1582 897 1593 931
rect 1520 885 1593 897
rect 1793 944 1929 969
rect 1793 910 1804 944
rect 1838 931 1929 944
rect 1838 910 1884 931
rect 1793 897 1884 910
rect 1918 897 1929 931
rect 1793 885 1929 897
rect 2029 1173 2082 1185
rect 2029 1139 2040 1173
rect 2074 1139 2082 1173
rect 2029 1093 2082 1139
rect 2029 1059 2040 1093
rect 2074 1059 2082 1093
rect 2029 1011 2082 1059
rect 2029 977 2040 1011
rect 2074 977 2082 1011
rect 2029 931 2082 977
rect 2029 897 2040 931
rect 2074 897 2082 931
rect 2029 885 2082 897
rect 1520 677 1578 689
rect 1520 643 1536 677
rect 1570 647 1578 677
rect 1808 677 1866 689
rect 1808 647 1816 677
rect 1570 643 1593 647
rect 626 607 679 619
rect 626 573 634 607
rect 668 573 679 607
rect 626 515 679 573
rect 626 481 634 515
rect 668 481 679 515
rect 626 469 679 481
rect 779 607 835 619
rect 779 573 790 607
rect 824 573 835 607
rect 779 515 835 573
rect 779 481 790 515
rect 824 481 835 515
rect 779 469 835 481
rect 935 607 988 619
rect 935 573 946 607
rect 980 573 988 607
rect 935 515 988 573
rect 1520 609 1593 643
rect 1520 575 1548 609
rect 1582 575 1593 609
rect 1520 563 1593 575
rect 1793 643 1816 647
rect 1850 643 1866 677
rect 1793 609 1866 643
rect 1793 575 1804 609
rect 1838 575 1866 609
rect 1793 563 1866 575
rect 935 481 946 515
rect 980 481 988 515
rect 935 469 988 481
<< mvndiffc >>
rect 702 1475 736 1509
rect 702 1395 736 1429
rect 702 1313 736 1347
rect 702 1233 736 1267
rect 858 1475 892 1509
rect 858 1395 892 1429
rect 858 1313 892 1347
rect 858 1233 892 1267
rect 1014 1475 1048 1509
rect 1014 1395 1048 1429
rect 1014 1313 1048 1347
rect 1014 1233 1048 1267
rect 1170 1475 1204 1509
rect 1170 1395 1204 1429
rect 1170 1313 1204 1347
rect 1170 1233 1204 1267
rect 1326 1475 1360 1509
rect 1326 1395 1360 1429
rect 1884 1475 1918 1509
rect 1884 1383 1918 1417
rect 2040 1475 2074 1509
rect 2040 1383 2074 1417
rect 1326 1313 1360 1347
rect 1326 1233 1360 1267
rect 1208 361 1242 395
rect 634 245 668 279
rect 634 153 668 187
rect 790 245 824 279
rect 790 153 824 187
rect 946 245 980 279
rect 946 153 980 187
rect 1208 281 1242 315
rect 1208 199 1242 233
rect 1208 119 1242 153
rect 1364 361 1398 395
rect 1364 281 1398 315
rect 1364 199 1398 233
rect 1364 119 1398 153
rect 1520 361 1554 395
rect 1520 281 1554 315
rect 1520 199 1554 233
rect 1520 119 1554 153
rect 1676 361 1710 395
rect 1676 281 1710 315
rect 1676 199 1710 233
rect 1676 119 1710 153
rect 1832 361 1866 395
rect 1832 281 1866 315
rect 1832 199 1866 233
rect 1832 119 1866 153
<< mvpdiffc >>
rect 1536 965 1570 999
rect 1884 1139 1918 1173
rect 1884 1059 1918 1093
rect 1884 977 1918 1011
rect 1548 897 1582 931
rect 1804 910 1838 944
rect 1884 897 1918 931
rect 2040 1139 2074 1173
rect 2040 1059 2074 1093
rect 2040 977 2074 1011
rect 2040 897 2074 931
rect 1536 643 1570 677
rect 634 573 668 607
rect 634 481 668 515
rect 790 573 824 607
rect 790 481 824 515
rect 946 573 980 607
rect 1548 575 1582 609
rect 1816 643 1850 677
rect 1804 575 1838 609
rect 946 481 980 515
<< mvpsubdiff >>
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1663 1645
rect 1697 1611 1759 1645
rect 1793 1611 1855 1645
rect 1889 1611 1951 1645
rect 1985 1611 2047 1645
rect 2081 1611 2112 1645
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 94 831
rect 1735 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2112 831
rect 626 789 988 797
rect 626 687 718 789
rect 956 687 988 789
rect 626 679 988 687
<< mvpsubdiffcont >>
rect 31 1611 65 1645
rect 127 1611 161 1645
rect 223 1611 257 1645
rect 319 1611 353 1645
rect 415 1611 449 1645
rect 511 1611 545 1645
rect 607 1611 641 1645
rect 703 1611 737 1645
rect 799 1611 833 1645
rect 895 1611 929 1645
rect 991 1611 1025 1645
rect 1087 1611 1121 1645
rect 1183 1611 1217 1645
rect 1279 1611 1313 1645
rect 1375 1611 1409 1645
rect 1471 1611 1505 1645
rect 1567 1611 1601 1645
rect 1663 1611 1697 1645
rect 1759 1611 1793 1645
rect 1855 1611 1889 1645
rect 1951 1611 1985 1645
rect 2047 1611 2081 1645
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 718 687 956 789
<< poly >>
rect 747 1521 847 1547
rect 903 1521 1003 1547
rect 1059 1521 1159 1547
rect 1215 1521 1315 1547
rect 1929 1521 2029 1547
rect 1929 1311 2029 1371
rect 1727 1295 2029 1311
rect 1727 1261 1743 1295
rect 1777 1261 2029 1295
rect 1727 1245 2029 1261
rect 1727 1227 1793 1245
rect 747 1199 847 1221
rect 903 1199 1003 1221
rect 1059 1199 1159 1221
rect 1215 1199 1315 1221
rect 747 1133 1315 1199
rect 1727 1193 1743 1227
rect 1777 1193 1793 1227
rect 1727 1159 1793 1193
rect 1929 1185 2029 1245
rect 930 1083 1132 1133
rect 930 1049 946 1083
rect 980 1049 1014 1083
rect 1048 1049 1082 1083
rect 1116 1049 1132 1083
rect 930 1033 1132 1049
rect 1727 1125 1743 1159
rect 1777 1125 1793 1159
rect 1727 1091 1793 1125
rect 1727 1057 1743 1091
rect 1777 1057 1793 1091
rect 1727 995 1793 1057
rect 1593 969 1793 995
rect 1593 859 1793 885
rect 1929 859 2029 885
rect 1475 771 1659 787
rect 1475 737 1491 771
rect 1525 737 1559 771
rect 1593 737 1659 771
rect 1475 721 1659 737
rect 679 619 779 645
rect 835 619 935 645
rect 1593 673 1659 721
rect 1593 647 1793 673
rect 1593 537 1793 563
rect 1112 479 1821 495
rect 499 424 565 440
rect 499 390 515 424
rect 549 407 565 424
rect 679 407 779 469
rect 549 390 779 407
rect 499 356 779 390
rect 499 322 515 356
rect 549 341 779 356
rect 549 322 565 341
rect 499 306 565 322
rect 679 291 779 341
rect 835 407 935 469
rect 1112 445 1128 479
rect 1162 445 1196 479
rect 1230 445 1264 479
rect 1298 445 1821 479
rect 1112 429 1821 445
rect 1253 407 1353 429
rect 1409 407 1509 429
rect 1565 407 1665 429
rect 1721 407 1821 429
rect 835 391 969 407
rect 835 357 851 391
rect 885 357 919 391
rect 953 357 969 391
rect 835 341 969 357
rect 835 291 935 341
rect 679 115 779 141
rect 835 115 935 141
rect 1253 81 1353 107
rect 1409 81 1509 107
rect 1565 81 1665 107
rect 1721 81 1821 107
<< polycont >>
rect 1743 1261 1777 1295
rect 1743 1193 1777 1227
rect 946 1049 980 1083
rect 1014 1049 1048 1083
rect 1082 1049 1116 1083
rect 1743 1125 1777 1159
rect 1743 1057 1777 1091
rect 1491 737 1525 771
rect 1559 737 1593 771
rect 515 390 549 424
rect 515 322 549 356
rect 1128 445 1162 479
rect 1196 445 1230 479
rect 1264 445 1298 479
rect 851 357 885 391
rect 919 357 953 391
<< locali >>
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1663 1645
rect 1697 1611 1759 1645
rect 1793 1611 1855 1645
rect 1889 1611 1951 1645
rect 1985 1611 2047 1645
rect 2081 1611 2112 1645
rect 660 1543 1402 1577
rect 660 1509 666 1543
rect 700 1509 738 1543
rect 772 1509 778 1543
rect 972 1509 978 1543
rect 1012 1509 1050 1543
rect 1084 1509 1090 1543
rect 1284 1509 1290 1543
rect 1324 1509 1362 1543
rect 1396 1509 1402 1543
rect 660 1475 702 1509
rect 736 1475 778 1509
rect 660 1429 778 1475
rect 660 1395 702 1429
rect 736 1395 778 1429
rect 660 1347 778 1395
rect 660 1313 702 1347
rect 736 1313 778 1347
rect 660 1267 778 1313
rect 660 1233 702 1267
rect 736 1233 778 1267
rect 660 1217 778 1233
rect 842 1475 858 1509
rect 892 1475 908 1509
rect 842 1429 908 1475
rect 842 1395 858 1429
rect 892 1395 908 1429
rect 842 1347 908 1395
rect 842 1313 858 1347
rect 892 1313 908 1347
rect 842 1267 908 1313
rect 842 1233 858 1267
rect 892 1233 908 1267
rect 972 1475 1014 1509
rect 1048 1475 1090 1509
rect 972 1429 1090 1475
rect 972 1395 1014 1429
rect 1048 1395 1090 1429
rect 972 1347 1090 1395
rect 972 1313 1014 1347
rect 1048 1313 1090 1347
rect 972 1267 1090 1313
rect 972 1233 1014 1267
rect 1048 1233 1090 1267
rect 1154 1475 1170 1509
rect 1204 1475 1220 1509
rect 1154 1429 1220 1475
rect 1154 1395 1170 1429
rect 1204 1395 1220 1429
rect 1154 1347 1220 1395
rect 1154 1313 1170 1347
rect 1204 1313 1220 1347
rect 1154 1267 1220 1313
rect 1154 1233 1170 1267
rect 1204 1233 1220 1267
rect 1284 1475 1326 1509
rect 1360 1475 1402 1509
rect 1284 1429 1402 1475
rect 1284 1395 1326 1429
rect 1360 1395 1402 1429
rect 1284 1347 1402 1395
rect 1842 1543 1960 1549
rect 1842 1509 1848 1543
rect 1882 1509 1920 1543
rect 1954 1509 1960 1543
rect 1842 1475 1884 1509
rect 1918 1475 1960 1509
rect 1842 1417 1960 1475
rect 1842 1383 1884 1417
rect 1918 1383 1960 1417
rect 1842 1367 1960 1383
rect 2024 1509 2090 1525
rect 2024 1475 2040 1509
rect 2074 1475 2090 1509
rect 2024 1417 2090 1475
rect 2024 1383 2040 1417
rect 2074 1383 2090 1417
rect 1284 1313 1326 1347
rect 1360 1313 1402 1347
rect 1284 1267 1402 1313
rect 1284 1233 1326 1267
rect 1360 1233 1402 1267
rect 1727 1295 1793 1311
rect 1727 1261 1743 1295
rect 1777 1261 1793 1295
rect 842 1199 908 1233
rect 1154 1199 1220 1233
rect 1727 1227 1793 1261
rect 842 1133 1586 1199
rect 618 1083 1132 1099
rect 618 1049 946 1083
rect 980 1049 1014 1083
rect 1048 1049 1082 1083
rect 1116 1049 1132 1083
rect 618 1033 1132 1049
rect 0 797 31 831
rect 65 797 160 831
rect 618 607 684 1033
rect 1520 999 1586 1133
rect 1727 1193 1743 1227
rect 1777 1193 1793 1227
rect 1727 1159 1793 1193
rect 1727 1125 1743 1159
rect 1777 1125 1793 1159
rect 1727 1107 1793 1125
rect 1520 965 1536 999
rect 1570 965 1586 999
rect 1520 931 1586 965
rect 1520 897 1548 931
rect 1582 897 1586 931
rect 718 789 956 805
rect 1520 787 1586 897
rect 1643 1091 1793 1107
rect 1643 1057 1743 1091
rect 1777 1057 1793 1091
rect 1643 1041 1793 1057
rect 1842 1173 1960 1189
rect 1842 1139 1884 1173
rect 1918 1139 1960 1173
rect 1842 1093 1960 1139
rect 1842 1059 1884 1093
rect 1918 1059 1960 1093
rect 1475 771 1609 787
rect 1475 737 1491 771
rect 1525 737 1559 771
rect 1593 737 1609 771
rect 1475 721 1609 737
rect 718 671 956 687
rect 1520 677 1586 687
rect 618 573 634 607
rect 668 573 684 607
rect 618 515 684 573
rect 618 481 634 515
rect 668 481 684 515
rect 499 424 561 440
rect 499 390 515 424
rect 549 390 561 424
rect 499 356 561 390
rect 499 322 515 356
rect 549 322 561 356
rect 499 306 561 322
rect 618 399 684 481
rect 748 644 866 671
rect 748 610 754 644
rect 788 610 826 644
rect 860 610 866 644
rect 1520 643 1536 677
rect 1570 643 1586 677
rect 1520 625 1586 643
rect 1643 625 1709 1041
rect 1842 1011 1960 1059
rect 1842 977 1884 1011
rect 1918 977 1960 1011
rect 1842 960 1960 977
rect 1758 944 1960 960
rect 1758 933 1804 944
rect 1838 933 1960 944
rect 1758 899 1776 933
rect 1838 910 1848 933
rect 1810 899 1848 910
rect 1882 931 1920 933
rect 1882 899 1884 931
rect 1758 897 1884 899
rect 1918 899 1920 931
rect 1954 899 1960 933
rect 1918 897 1960 899
rect 1758 881 1960 897
rect 2024 1173 2090 1383
rect 2024 1139 2040 1173
rect 2074 1139 2090 1173
rect 2024 1093 2090 1139
rect 2024 1059 2040 1093
rect 2074 1059 2090 1093
rect 2024 1011 2090 1059
rect 2024 977 2040 1011
rect 2074 977 2090 1011
rect 2024 931 2090 977
rect 2024 897 2040 931
rect 2074 897 2090 931
rect 2024 881 2090 897
rect 1743 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2112 831
rect 748 607 866 610
rect 748 573 790 607
rect 824 573 866 607
rect 748 515 866 573
rect 748 481 790 515
rect 824 481 866 515
rect 748 465 866 481
rect 930 607 996 623
rect 930 573 946 607
rect 980 573 996 607
rect 930 515 996 573
rect 1520 609 1709 625
rect 1520 575 1548 609
rect 1582 575 1709 609
rect 1520 559 1709 575
rect 1788 729 1906 741
rect 1788 695 1794 729
rect 1828 695 1866 729
rect 1900 695 1906 729
rect 1788 677 1906 695
rect 1788 643 1816 677
rect 1850 643 1906 677
rect 1788 609 1906 643
rect 1788 575 1804 609
rect 1838 575 1906 609
rect 1788 559 1906 575
rect 930 481 946 515
rect 980 495 996 515
rect 1643 495 1709 559
rect 980 481 1314 495
rect 930 479 1314 481
rect 930 445 1128 479
rect 1162 445 1196 479
rect 1230 445 1264 479
rect 1298 445 1314 479
rect 930 433 1314 445
rect 1066 429 1314 433
rect 1348 429 1726 495
rect 618 391 969 399
rect 618 357 851 391
rect 885 357 919 391
rect 953 357 969 391
rect 618 349 969 357
rect 618 279 684 349
rect 1066 295 1132 429
rect 1348 395 1414 429
rect 1660 395 1726 429
rect 618 245 634 279
rect 668 245 684 279
rect 618 187 684 245
rect 618 153 634 187
rect 668 153 684 187
rect 618 137 684 153
rect 748 279 866 295
rect 748 245 790 279
rect 824 245 866 279
rect 748 187 866 245
rect 748 153 790 187
rect 824 153 866 187
rect 748 119 866 153
rect 930 279 1132 295
rect 930 245 946 279
rect 980 245 1132 279
rect 930 229 1132 245
rect 1166 361 1208 395
rect 1242 361 1284 395
rect 1166 315 1284 361
rect 1166 281 1208 315
rect 1242 281 1284 315
rect 1166 233 1284 281
rect 930 187 996 229
rect 930 153 946 187
rect 980 153 996 187
rect 930 137 996 153
rect 1166 199 1208 233
rect 1242 199 1284 233
rect 1166 153 1284 199
rect 748 85 754 119
rect 788 85 826 119
rect 860 85 866 119
rect 1166 119 1208 153
rect 1242 119 1284 153
rect 1348 361 1364 395
rect 1398 361 1414 395
rect 1348 315 1414 361
rect 1348 281 1364 315
rect 1398 281 1414 315
rect 1348 233 1414 281
rect 1348 199 1364 233
rect 1398 199 1414 233
rect 1348 153 1414 199
rect 1348 119 1364 153
rect 1398 119 1414 153
rect 1478 361 1520 395
rect 1554 361 1596 395
rect 1478 315 1596 361
rect 1478 281 1520 315
rect 1554 281 1596 315
rect 1478 233 1596 281
rect 1478 199 1520 233
rect 1554 199 1596 233
rect 1478 153 1596 199
rect 1478 119 1520 153
rect 1554 119 1596 153
rect 1660 361 1676 395
rect 1710 361 1726 395
rect 1660 315 1726 361
rect 1660 281 1676 315
rect 1710 281 1726 315
rect 1660 233 1726 281
rect 1660 199 1676 233
rect 1710 199 1726 233
rect 1660 153 1726 199
rect 1660 119 1676 153
rect 1710 119 1726 153
rect 1790 361 1832 395
rect 1866 361 1908 395
rect 1790 315 1908 361
rect 1790 281 1832 315
rect 1866 281 1908 315
rect 1790 233 1908 281
rect 1790 199 1832 233
rect 1866 199 1908 233
rect 1790 153 1908 199
rect 1790 119 1832 153
rect 1866 119 1908 153
rect 1166 85 1172 119
rect 1206 85 1244 119
rect 1278 85 1284 119
rect 1478 85 1484 119
rect 1518 85 1556 119
rect 1590 85 1596 119
rect 1790 85 1796 119
rect 1830 85 1868 119
rect 1902 85 1908 119
rect 748 51 1908 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< viali >>
rect 31 1611 65 1645
rect 127 1611 161 1645
rect 223 1611 257 1645
rect 319 1611 353 1645
rect 415 1611 449 1645
rect 511 1611 545 1645
rect 607 1611 641 1645
rect 703 1611 737 1645
rect 799 1611 833 1645
rect 895 1611 929 1645
rect 991 1611 1025 1645
rect 1087 1611 1121 1645
rect 1183 1611 1217 1645
rect 1279 1611 1313 1645
rect 1375 1611 1409 1645
rect 1471 1611 1505 1645
rect 1567 1611 1601 1645
rect 1663 1611 1697 1645
rect 1759 1611 1793 1645
rect 1855 1611 1889 1645
rect 1951 1611 1985 1645
rect 2047 1611 2081 1645
rect 666 1509 700 1543
rect 738 1509 772 1543
rect 978 1509 1012 1543
rect 1050 1509 1084 1543
rect 1290 1509 1324 1543
rect 1362 1509 1396 1543
rect 1848 1509 1882 1543
rect 1920 1509 1954 1543
rect 31 797 65 831
rect 754 610 788 644
rect 826 610 860 644
rect 1776 910 1804 933
rect 1804 910 1810 933
rect 1776 899 1810 910
rect 1848 899 1882 933
rect 1920 899 1954 933
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 1794 695 1828 729
rect 1866 695 1900 729
rect 754 85 788 119
rect 826 85 860 119
rect 1172 85 1206 119
rect 1244 85 1278 119
rect 1484 85 1518 119
rect 1556 85 1590 119
rect 1796 85 1830 119
rect 1868 85 1902 119
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 1645 2112 1651
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1663 1645
rect 1697 1611 1759 1645
rect 1793 1611 1855 1645
rect 1889 1611 1951 1645
rect 1985 1611 2047 1645
rect 2081 1611 2112 1645
rect 0 1605 2112 1611
rect 0 1543 2112 1577
rect 0 1509 666 1543
rect 700 1509 738 1543
rect 772 1509 978 1543
rect 1012 1509 1050 1543
rect 1084 1509 1290 1543
rect 1324 1509 1362 1543
rect 1396 1509 1848 1543
rect 1882 1509 1920 1543
rect 1954 1509 2112 1543
rect 0 1503 2112 1509
rect 0 933 2112 939
rect 0 899 1776 933
rect 1810 899 1848 933
rect 1882 899 1920 933
rect 1954 899 2112 933
rect 0 865 2112 899
rect 0 831 2112 837
rect 0 797 31 831
rect 65 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2112 831
rect 0 791 2112 797
rect 0 729 2112 763
rect 0 695 1794 729
rect 1828 695 1866 729
rect 1900 695 2112 729
rect 0 689 2112 695
rect 14 644 2098 661
rect 14 610 754 644
rect 788 610 826 644
rect 860 610 2098 644
rect 14 604 2098 610
rect 0 119 2112 125
rect 0 85 754 119
rect 788 85 826 119
rect 860 85 1172 119
rect 1206 85 1244 119
rect 1278 85 1484 119
rect 1518 85 1556 119
rect 1590 85 1796 119
rect 1830 85 1868 119
rect 1902 85 2112 119
rect 0 51 2112 85
rect 0 17 2112 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -23 2112 -17
<< labels >>
rlabel comment s 0 0 0 0 4 lsbufhv2hv_lh_1
flabel metal1 s 0 865 2112 939 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 689 2112 763 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 1503 2112 1577 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 51 2112 125 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 0 2112 23 0 FreeSans 340 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 14 604 2098 661 0 FreeSans 340 0 0 0 LOWHVPWR
port 2 nsew power bidirectional
flabel metal1 s 0 791 2112 837 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 0 1605 2112 1628 0 FreeSans 340 0 0 0 VNB
port 4 nsew ground bidirectional
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 2047 1204 2081 1238 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 2047 1130 2081 1164 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 2047 1056 2081 1090 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 2047 1278 2081 1312 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 2047 1352 2081 1386 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
rlabel viali s 826 610 860 644 1 LOWHVPWR
port 2 nsew power bidirectional
rlabel viali s 754 610 788 644 1 LOWHVPWR
port 2 nsew power bidirectional
rlabel metal1 s 14 604 2098 661 1 LOWHVPWR
port 2 nsew power bidirectional
rlabel locali s 1790 85 1908 395 1 VGND
port 3 nsew ground bidirectional
rlabel locali s 1478 85 1596 395 1 VGND
port 3 nsew ground bidirectional
rlabel locali s 1166 85 1284 395 1 VGND
port 3 nsew ground bidirectional
rlabel locali s 748 85 866 295 1 VGND
port 3 nsew ground bidirectional
rlabel locali s 748 51 1908 85 1 VGND
port 3 nsew ground bidirectional
rlabel locali s 1842 1367 1960 1549 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 1920 1509 1954 1543 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 1868 85 1902 119 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 1848 1509 1882 1543 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 1796 85 1830 119 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 1556 85 1590 119 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 1484 85 1518 119 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 1362 1509 1396 1543 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 1290 1509 1324 1543 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 1244 85 1278 119 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 1172 85 1206 119 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 1050 1509 1084 1543 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 978 1509 1012 1543 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 826 85 860 119 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 754 85 788 119 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 738 1509 772 1543 1 VGND
port 3 nsew ground bidirectional
rlabel viali s 666 1509 700 1543 1 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 51 2112 125 1 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 1503 2112 1577 1 VGND
port 3 nsew ground bidirectional
rlabel locali s 0 1611 2112 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 2047 1611 2081 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 2047 -17 2081 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1951 1611 1985 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1951 -17 1985 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1855 1611 1889 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1855 -17 1889 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1759 1611 1793 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1759 -17 1793 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1663 1611 1697 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1663 -17 1697 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1567 1611 1601 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1567 -17 1601 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1471 1611 1505 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1471 -17 1505 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1375 1611 1409 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1375 -17 1409 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1279 1611 1313 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1279 -17 1313 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1183 1611 1217 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1183 -17 1217 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1087 1611 1121 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 1087 -17 1121 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 991 1611 1025 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 991 -17 1025 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 895 1611 929 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 895 -17 929 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 799 1611 833 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 799 -17 833 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 703 1611 737 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 703 -17 737 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 607 1611 641 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 607 -17 641 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 511 1611 545 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 511 -17 545 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 415 1611 449 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 415 -17 449 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 319 1611 353 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 319 -17 353 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 223 1611 257 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 223 -17 257 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 127 1611 161 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 127 -17 161 17 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 31 1611 65 1645 1 VNB
port 4 nsew ground bidirectional
rlabel viali s 31 -17 65 17 1 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 -23 2112 23 1 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 1605 2112 1651 1 VNB
port 4 nsew ground bidirectional
rlabel locali s 1743 797 2112 831 1 VPB
port 5 nsew power bidirectional
rlabel viali s 2047 797 2081 831 1 VPB
port 5 nsew power bidirectional
rlabel viali s 1951 797 1985 831 1 VPB
port 5 nsew power bidirectional
rlabel viali s 1855 797 1889 831 1 VPB
port 5 nsew power bidirectional
rlabel viali s 1759 797 1793 831 1 VPB
port 5 nsew power bidirectional
rlabel viali s 31 797 65 831 1 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 791 2112 837 1 VPB
port 5 nsew power bidirectional
rlabel locali s 1788 559 1906 741 1 VPWR
port 6 nsew power bidirectional
rlabel viali s 1920 899 1954 933 1 VPWR
port 6 nsew power bidirectional
rlabel viali s 1866 695 1900 729 1 VPWR
port 6 nsew power bidirectional
rlabel viali s 1848 899 1882 933 1 VPWR
port 6 nsew power bidirectional
rlabel viali s 1794 695 1828 729 1 VPWR
port 6 nsew power bidirectional
rlabel viali s 1776 899 1810 933 1 VPWR
port 6 nsew power bidirectional
rlabel metal1 s 0 689 2112 763 1 VPWR
port 6 nsew power bidirectional
rlabel metal1 s 0 865 2112 939 1 VPWR
port 6 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 2112 1628
string GDS_END 167916
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 146448
string LEFclass CORE
string LEFsite unithvdbl
string LEFsymmetry X Y
<< end >>
