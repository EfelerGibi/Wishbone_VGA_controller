magic
tech sky130A
magscale 1 2
timestamp 1683767628
use sky130_fd_pr__hvdfm1sd2__example_5595914180829  sky130_fd_pr__hvdfm1sd2__example_5595914180829_0
timestamp 1683767628
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180829  sky130_fd_pr__hvdfm1sd2__example_5595914180829_1
timestamp 1683767628
transform 1 0 180 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 27758142
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 27757152
<< end >>
