magic
tech sky130A
timestamp 1683767628
<< properties >>
string GDS_END 7197292
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7196588
<< end >>
