magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< metal4 >>
rect 0 41065 1000 45908
rect 0 19915 1000 24908
rect 0 18725 1000 19615
rect 0 17555 1000 18445
rect 0 17189 1000 17255
rect 0 16533 1000 17129
rect 0 16237 48 16473
rect 284 16237 380 16473
rect 616 16237 711 16473
rect 947 16237 1000 16473
rect 0 15581 1000 16177
rect 0 15455 1000 15521
rect 0 14225 1000 15155
rect 0 13255 1000 13945
rect 0 12285 1000 12975
rect 0 11075 1000 12005
rect 0 9865 1000 10795
rect 0 8895 1000 9585
rect 0 7685 1000 8615
rect 0 6315 1000 7405
<< via4 >>
rect 48 16237 284 16473
rect 380 16237 616 16473
rect 711 16237 947 16473
<< metal5 >>
rect 0 41065 1000 45908
rect 0 19915 1000 24905
rect 0 18745 1000 19595
rect 0 17575 1000 18425
rect 0 16473 1000 17255
rect 0 16237 48 16473
rect 284 16237 380 16473
rect 616 16237 711 16473
rect 947 16237 1000 16473
rect 0 15455 1000 16237
rect 0 14245 1000 15135
rect 0 13275 1000 13925
rect 0 12305 1000 12955
rect 0 11095 1000 11985
rect 0 9885 1000 10775
rect 0 8915 1000 9565
rect 0 7705 1000 8595
rect 0 6335 1000 7385
<< properties >>
string GDS_END 194548
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 192176
<< end >>
