magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 157 186 203
rect 1 21 735 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 175 47 205 131
rect 268 47 298 131
rect 459 47 489 131
rect 543 47 573 131
rect 627 47 657 131
<< scpmoshvt >>
rect 79 297 109 497
rect 176 369 206 453
rect 286 369 316 453
rect 461 369 491 453
rect 555 369 585 453
rect 627 369 657 453
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 131 160 177
rect 109 122 175 131
rect 109 88 124 122
rect 158 88 175 122
rect 109 47 175 88
rect 205 47 268 131
rect 298 113 350 131
rect 298 79 308 113
rect 342 79 350 113
rect 298 47 350 79
rect 407 114 459 131
rect 407 80 415 114
rect 449 80 459 114
rect 407 47 459 80
rect 489 114 543 131
rect 489 80 499 114
rect 533 80 543 114
rect 489 47 543 80
rect 573 95 627 131
rect 573 61 583 95
rect 617 61 627 95
rect 573 47 627 61
rect 657 104 709 131
rect 657 70 667 104
rect 701 70 709 104
rect 657 47 709 70
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 297 79 375
rect 109 481 161 497
rect 109 447 119 481
rect 153 453 161 481
rect 332 481 446 493
rect 332 453 366 481
rect 153 447 176 453
rect 109 369 176 447
rect 206 369 286 453
rect 316 447 366 453
rect 400 453 446 481
rect 400 447 461 453
rect 316 369 461 447
rect 491 429 555 453
rect 491 395 501 429
rect 535 395 555 429
rect 491 369 555 395
rect 585 369 627 453
rect 657 429 709 453
rect 657 395 667 429
rect 701 395 709 429
rect 657 369 709 395
rect 109 297 161 369
rect 221 343 271 369
rect 221 309 229 343
rect 263 309 271 343
rect 221 297 271 309
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 124 88 158 122
rect 308 79 342 113
rect 415 80 449 114
rect 499 80 533 114
rect 583 61 617 95
rect 667 70 701 104
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 447 153 481
rect 366 447 400 481
rect 501 395 535 429
rect 667 395 701 429
rect 229 309 263 343
<< poly >>
rect 79 497 109 523
rect 176 453 206 479
rect 286 453 316 479
rect 461 453 491 479
rect 555 453 585 479
rect 627 453 657 479
rect 79 265 109 297
rect 176 265 206 369
rect 76 249 130 265
rect 76 215 86 249
rect 120 215 130 249
rect 76 199 130 215
rect 172 249 226 265
rect 172 215 182 249
rect 216 215 226 249
rect 286 220 316 369
rect 461 337 491 369
rect 358 321 491 337
rect 358 287 368 321
rect 402 312 491 321
rect 402 287 489 312
rect 358 271 489 287
rect 172 199 226 215
rect 268 204 326 220
rect 79 177 109 199
rect 175 131 205 199
rect 268 170 278 204
rect 312 170 326 204
rect 268 154 326 170
rect 268 131 298 154
rect 459 131 489 271
rect 555 265 585 369
rect 531 249 585 265
rect 531 215 541 249
rect 575 215 585 249
rect 531 199 585 215
rect 627 265 657 369
rect 627 249 715 265
rect 627 215 666 249
rect 700 215 715 249
rect 627 199 715 215
rect 543 131 573 199
rect 627 131 657 199
rect 79 21 109 47
rect 175 21 205 47
rect 268 21 298 47
rect 459 21 489 47
rect 543 21 573 47
rect 627 21 657 47
<< polycont >>
rect 86 215 120 249
rect 182 215 216 249
rect 368 287 402 321
rect 278 170 312 204
rect 541 215 575 249
rect 666 215 700 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 477 69 493
rect 17 443 35 477
rect 103 481 169 527
rect 103 447 119 481
rect 153 447 169 481
rect 343 481 423 527
rect 343 447 366 481
rect 400 447 423 481
rect 17 409 69 443
rect 481 429 547 458
rect 481 411 501 429
rect 17 375 35 409
rect 17 359 69 375
rect 131 395 501 411
rect 535 395 547 429
rect 131 377 547 395
rect 17 165 52 359
rect 131 323 165 377
rect 86 289 165 323
rect 199 309 229 343
rect 263 321 402 343
rect 263 309 368 321
rect 199 299 368 309
rect 86 249 120 289
rect 347 287 368 299
rect 347 271 402 287
rect 436 299 547 377
rect 154 249 244 255
rect 154 215 182 249
rect 216 215 244 249
rect 86 199 120 215
rect 278 204 313 220
rect 214 170 278 181
rect 312 170 313 204
rect 17 161 85 165
rect 17 127 35 161
rect 69 127 85 161
rect 17 93 85 127
rect 17 59 35 93
rect 69 59 85 93
rect 17 51 85 59
rect 124 122 158 150
rect 124 17 158 88
rect 214 147 313 170
rect 214 76 258 147
rect 347 113 381 271
rect 436 249 470 299
rect 581 265 616 485
rect 650 429 719 527
rect 650 395 667 429
rect 701 395 719 429
rect 650 363 719 395
rect 431 215 470 249
rect 504 249 616 265
rect 504 215 541 249
rect 575 215 616 249
rect 650 249 719 329
rect 650 215 666 249
rect 700 215 719 249
rect 431 138 465 215
rect 292 79 308 113
rect 342 79 381 113
rect 415 114 465 138
rect 449 80 465 114
rect 415 64 465 80
rect 499 145 719 181
rect 499 114 549 145
rect 533 80 549 114
rect 499 64 549 80
rect 583 95 617 111
rect 651 104 719 145
rect 651 70 667 104
rect 701 70 719 104
rect 651 64 719 70
rect 583 17 617 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 210 221 244 255 0 FreeSans 400 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 30 425 64 459 0 FreeSans 400 0 0 0 X
port 9 nsew signal output
flabel locali s 214 85 248 119 0 FreeSans 400 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 581 289 615 323 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel locali s 673 221 707 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 o2bb2a_1
rlabel metal1 s 0 -48 736 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 1216942
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1210550
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 3.680 0.000 
<< end >>
