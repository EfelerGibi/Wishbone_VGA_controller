magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 1 21 1239 203
rect 30 -17 64 21
<< locali >>
rect 919 391 953 493
rect 1087 391 1121 493
rect 907 357 1259 391
rect 30 289 571 323
rect 30 215 105 289
rect 145 215 211 249
rect 271 215 341 255
rect 397 215 463 255
rect 505 215 571 289
rect 161 181 195 215
rect 397 181 434 215
rect 161 147 434 181
rect 715 215 806 257
rect 763 149 806 215
rect 1225 165 1259 357
rect 901 131 1259 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 35 391 69 493
rect 103 425 169 527
rect 203 391 237 493
rect 271 425 337 527
rect 371 391 405 493
rect 439 425 505 527
rect 563 459 765 493
rect 563 391 597 459
rect 35 357 597 391
rect 631 325 697 423
rect 731 359 765 459
rect 819 425 885 527
rect 987 425 1053 527
rect 1155 425 1221 527
rect 631 291 879 325
rect 35 17 69 181
rect 631 174 669 291
rect 845 265 879 291
rect 470 161 669 174
rect 470 140 697 161
rect 845 199 1187 265
rect 470 113 504 140
rect 271 79 504 113
rect 540 17 597 106
rect 631 59 697 140
rect 747 17 853 113
rect 987 17 1053 97
rect 1155 17 1221 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
rlabel locali s 271 215 341 255 6 A1
port 1 nsew signal input
rlabel locali s 161 147 434 181 6 A2
port 2 nsew signal input
rlabel locali s 397 181 434 215 6 A2
port 2 nsew signal input
rlabel locali s 161 181 195 215 6 A2
port 2 nsew signal input
rlabel locali s 397 215 463 255 6 A2
port 2 nsew signal input
rlabel locali s 145 215 211 249 6 A2
port 2 nsew signal input
rlabel locali s 505 215 571 289 6 A3
port 3 nsew signal input
rlabel locali s 30 215 105 289 6 A3
port 3 nsew signal input
rlabel locali s 30 289 571 323 6 A3
port 3 nsew signal input
rlabel locali s 763 149 806 215 6 B1
port 4 nsew signal input
rlabel locali s 715 215 806 257 6 B1
port 4 nsew signal input
rlabel metal1 s 0 -48 1288 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 1239 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1326 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1288 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 901 131 1259 165 6 X
port 9 nsew signal output
rlabel locali s 1225 165 1259 357 6 X
port 9 nsew signal output
rlabel locali s 907 357 1259 391 6 X
port 9 nsew signal output
rlabel locali s 1087 391 1121 493 6 X
port 9 nsew signal output
rlabel locali s 919 391 953 493 6 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1288 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 4137538
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4127676
<< end >>
