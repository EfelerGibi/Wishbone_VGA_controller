magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< locali >>
rect 0 1396 2554 1432
rect 1856 902 1890 918
rect 1855 868 1856 885
rect 1855 852 1890 868
rect 1855 724 1889 852
rect 1558 698 1592 714
rect 1855 698 2051 724
rect 1694 690 2051 698
rect 2276 690 2395 724
rect 1694 664 1889 690
rect 1558 648 1592 664
rect 2361 520 2395 690
rect 2361 470 2395 486
rect 0 -18 2554 18
<< viali >>
rect 1856 868 1890 902
rect 1558 664 1592 698
rect 2361 486 2395 520
<< metal1 >>
rect 1840 859 1846 911
rect 1898 859 1905 911
rect 1543 655 1549 707
rect 1601 655 1607 707
rect 2346 477 2352 529
rect 2404 477 2410 529
<< via1 >>
rect 1846 902 1898 911
rect 1846 868 1856 902
rect 1856 868 1890 902
rect 1890 868 1898 902
rect 1846 859 1898 868
rect 1549 698 1601 707
rect 1549 664 1558 698
rect 1558 664 1592 698
rect 1592 664 1601 698
rect 1549 655 1601 664
rect 2352 520 2404 529
rect 2352 486 2361 520
rect 2361 486 2395 520
rect 2395 486 2404 520
rect 2352 477 2404 486
<< metal2 >>
rect 1846 911 1898 917
rect 1846 853 1898 859
rect 369 692 423 756
rect 1549 707 1601 713
rect 1115 655 1549 661
rect 1115 609 1601 655
rect 137 538 203 590
rect 2352 529 2404 535
rect 2352 471 2404 477
use sky130_fd_bd_sram__openram_dff_2  sky130_fd_bd_sram__openram_dff_0
timestamp 1683767628
transform 1 0 0 0 1 0
box -36 -43 1204 1467
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_0
timestamp 1683767628
transform 1 0 1844 0 1 852
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1
timestamp 1683767628
transform 1 0 2349 0 1 470
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_2
timestamp 1683767628
transform 1 0 1546 0 1 648
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_0
timestamp 1683767628
transform 1 0 1840 0 1 853
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_1
timestamp 1683767628
transform 1 0 2346 0 1 471
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_2
timestamp 1683767628
transform 1 0 1543 0 1 649
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_pinv_2  sky130_sram_2kbyte_1rw1r_32x512_8_pinv_2_0
timestamp 1683767628
transform 1 0 1494 0 1 0
box -36 -17 512 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_pinv_3  sky130_sram_2kbyte_1rw1r_32x512_8_pinv_3_0
timestamp 1683767628
transform 1 0 1970 0 1 0
box -36 -17 620 1471
<< labels >>
rlabel metal2 s 369 692 423 756 4 clk
port 1 nsew
rlabel metal2 s 137 538 203 590 4 D
port 2 nsew
rlabel metal2 s 2364 489 2392 517 4 Q
port 3 nsew
rlabel metal2 s 1858 871 1886 899 4 Qb
port 4 nsew
rlabel locali s 1277 1414 1277 1414 4 vdd
rlabel locali s 1277 0 1277 0 4 gnd
<< properties >>
string FIXED_BBOX 0 0 2554 1414
string GDS_END 395128
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 392482
<< end >>
