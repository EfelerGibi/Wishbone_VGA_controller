magic
tech sky130B
timestamp 1683767628
<< obsli1 >>
rect 0 1136 5573 1169
rect 0 33 14 1122
rect 28 47 42 1136
rect 56 33 70 1122
rect 84 47 98 1136
rect 112 33 126 1122
rect 140 47 154 1136
rect 168 33 182 1122
rect 196 47 210 1136
rect 224 33 238 1122
rect 252 47 266 1136
rect 280 33 294 1122
rect 308 47 322 1136
rect 336 33 350 1122
rect 364 47 378 1136
rect 392 33 406 1122
rect 420 47 434 1136
rect 448 33 462 1122
rect 476 47 490 1136
rect 504 33 518 1122
rect 532 47 546 1136
rect 560 33 574 1122
rect 588 47 602 1136
rect 616 33 630 1122
rect 644 47 658 1136
rect 672 33 686 1122
rect 700 47 714 1136
rect 728 33 742 1122
rect 756 47 770 1136
rect 784 33 798 1122
rect 812 47 826 1136
rect 840 33 854 1122
rect 868 47 882 1136
rect 896 33 910 1122
rect 924 47 938 1136
rect 952 33 966 1122
rect 980 47 994 1136
rect 1008 33 1022 1122
rect 1036 47 1050 1136
rect 1064 33 1078 1122
rect 1092 47 1106 1136
rect 1120 33 1134 1122
rect 1148 47 1162 1136
rect 1176 33 1190 1122
rect 1204 47 1218 1136
rect 1232 33 1246 1122
rect 1260 47 1274 1136
rect 1288 33 1302 1122
rect 1316 47 1330 1136
rect 1344 33 1358 1122
rect 1372 47 1386 1136
rect 1400 33 1414 1122
rect 1428 47 1442 1136
rect 1456 33 1470 1122
rect 1484 47 1498 1136
rect 1512 33 1526 1122
rect 1540 47 1554 1136
rect 1568 33 1582 1122
rect 1596 47 1610 1136
rect 1624 33 1638 1122
rect 1652 47 1666 1136
rect 1680 33 1694 1122
rect 1708 47 1722 1136
rect 1736 33 1750 1122
rect 1764 47 1778 1136
rect 1792 33 1806 1122
rect 1820 47 1834 1136
rect 1848 33 1862 1122
rect 1876 47 1890 1136
rect 1904 33 1918 1122
rect 1932 47 1946 1136
rect 1960 33 1974 1122
rect 1988 47 2002 1136
rect 2016 33 2030 1122
rect 2044 47 2058 1136
rect 2072 33 2086 1122
rect 2100 47 2114 1136
rect 2128 33 2142 1122
rect 2156 47 2170 1136
rect 2184 33 2198 1122
rect 2212 47 2226 1136
rect 2240 33 2254 1122
rect 2268 47 2282 1136
rect 2296 33 2310 1122
rect 2324 47 2338 1136
rect 2352 33 2366 1122
rect 2380 47 2394 1136
rect 2408 33 2422 1122
rect 2436 47 2450 1136
rect 2464 33 2478 1122
rect 2492 47 2506 1136
rect 2520 33 2534 1122
rect 2548 47 2562 1136
rect 2576 33 2590 1122
rect 2604 47 2618 1136
rect 2632 33 2646 1122
rect 2660 47 2674 1136
rect 2688 33 2702 1122
rect 2716 47 2730 1136
rect 2744 33 2758 1122
rect 2772 47 2786 1136
rect 2800 33 2814 1122
rect 2828 47 2842 1136
rect 2856 33 2870 1122
rect 2884 47 2898 1136
rect 2912 33 2926 1122
rect 2940 47 2954 1136
rect 2968 33 2982 1122
rect 2996 47 3010 1136
rect 3024 33 3038 1122
rect 3052 47 3066 1136
rect 3080 33 3094 1122
rect 3108 47 3122 1136
rect 3136 33 3150 1122
rect 3164 47 3178 1136
rect 3192 33 3206 1122
rect 3220 47 3234 1136
rect 3248 33 3262 1122
rect 3276 47 3290 1136
rect 3304 33 3318 1122
rect 3332 47 3346 1136
rect 3360 33 3374 1122
rect 3388 47 3402 1136
rect 3416 33 3430 1122
rect 3444 47 3458 1136
rect 3472 33 3486 1122
rect 3500 47 3514 1136
rect 3528 33 3542 1122
rect 3556 47 3570 1136
rect 3584 33 3598 1122
rect 3612 47 3626 1136
rect 3640 33 3654 1122
rect 3668 47 3682 1136
rect 3696 33 3710 1122
rect 3724 47 3738 1136
rect 3752 33 3766 1122
rect 3780 47 3794 1136
rect 3808 33 3822 1122
rect 3836 47 3850 1136
rect 3864 33 3878 1122
rect 3892 47 3906 1136
rect 3920 33 3934 1122
rect 3948 47 3962 1136
rect 3976 33 3990 1122
rect 4004 47 4018 1136
rect 4032 33 4046 1122
rect 4060 47 4074 1136
rect 4088 33 4102 1122
rect 4116 47 4130 1136
rect 4144 33 4158 1122
rect 4172 47 4186 1136
rect 4200 33 4214 1122
rect 4228 47 4242 1136
rect 4256 33 4270 1122
rect 4284 47 4298 1136
rect 4312 33 4326 1122
rect 4340 47 4354 1136
rect 4368 33 4382 1122
rect 4396 47 4410 1136
rect 4424 33 4438 1122
rect 4452 47 4466 1136
rect 4480 33 4494 1122
rect 4508 47 4522 1136
rect 4536 33 4550 1122
rect 4564 47 4578 1136
rect 4592 33 4606 1122
rect 4620 47 4634 1136
rect 4648 33 4662 1122
rect 4676 47 4690 1136
rect 4704 33 4718 1122
rect 4732 47 4746 1136
rect 4760 33 4774 1122
rect 4788 47 4802 1136
rect 4816 33 4830 1122
rect 4844 47 4858 1136
rect 4872 33 4886 1122
rect 4900 47 4914 1136
rect 4928 33 4942 1122
rect 4956 47 4970 1136
rect 4984 33 4998 1122
rect 5012 47 5026 1136
rect 5040 33 5054 1122
rect 5068 47 5082 1136
rect 5096 33 5110 1122
rect 5124 47 5138 1136
rect 5152 33 5166 1122
rect 5180 47 5194 1136
rect 5208 33 5222 1122
rect 5236 47 5250 1136
rect 5264 33 5278 1122
rect 5292 47 5306 1136
rect 5320 33 5334 1122
rect 5348 47 5362 1136
rect 5376 33 5390 1122
rect 5404 47 5418 1136
rect 5432 33 5446 1122
rect 5460 47 5474 1136
rect 5488 33 5502 1122
rect 5516 47 5530 1136
rect 5544 33 5573 1122
rect 0 0 5573 33
<< obsm1 >>
rect 0 1136 5573 1169
rect 0 47 14 1136
rect 28 33 42 1122
rect 56 47 70 1136
rect 84 33 98 1122
rect 112 47 126 1136
rect 140 33 154 1122
rect 168 47 182 1136
rect 196 33 210 1122
rect 224 47 238 1136
rect 252 33 266 1122
rect 280 47 294 1136
rect 308 33 322 1122
rect 336 47 350 1136
rect 364 33 378 1122
rect 392 47 406 1136
rect 420 33 434 1122
rect 448 47 462 1136
rect 476 33 490 1122
rect 504 47 518 1136
rect 532 33 546 1122
rect 560 47 574 1136
rect 588 33 602 1122
rect 616 47 630 1136
rect 644 33 658 1122
rect 672 47 686 1136
rect 700 33 714 1122
rect 728 47 742 1136
rect 756 33 770 1122
rect 784 47 798 1136
rect 812 33 826 1122
rect 840 47 854 1136
rect 868 33 882 1122
rect 896 47 910 1136
rect 924 33 938 1122
rect 952 47 966 1136
rect 980 33 994 1122
rect 1008 47 1022 1136
rect 1036 33 1050 1122
rect 1064 47 1078 1136
rect 1092 33 1106 1122
rect 1120 47 1134 1136
rect 1148 33 1162 1122
rect 1176 47 1190 1136
rect 1204 33 1218 1122
rect 1232 47 1246 1136
rect 1260 33 1274 1122
rect 1288 47 1302 1136
rect 1316 33 1330 1122
rect 1344 47 1358 1136
rect 1372 33 1386 1122
rect 1400 47 1414 1136
rect 1428 33 1442 1122
rect 1456 47 1470 1136
rect 1484 33 1498 1122
rect 1512 47 1526 1136
rect 1540 33 1554 1122
rect 1568 47 1582 1136
rect 1596 33 1610 1122
rect 1624 47 1638 1136
rect 1652 33 1666 1122
rect 1680 47 1694 1136
rect 1708 33 1722 1122
rect 1736 47 1750 1136
rect 1764 33 1778 1122
rect 1792 47 1806 1136
rect 1820 33 1834 1122
rect 1848 47 1862 1136
rect 1876 33 1890 1122
rect 1904 47 1918 1136
rect 1932 33 1946 1122
rect 1960 47 1974 1136
rect 1988 33 2002 1122
rect 2016 47 2030 1136
rect 2044 33 2058 1122
rect 2072 47 2086 1136
rect 2100 33 2114 1122
rect 2128 47 2142 1136
rect 2156 33 2170 1122
rect 2184 47 2198 1136
rect 2212 33 2226 1122
rect 2240 47 2254 1136
rect 2268 33 2282 1122
rect 2296 47 2310 1136
rect 2324 33 2338 1122
rect 2352 47 2366 1136
rect 2380 33 2394 1122
rect 2408 47 2422 1136
rect 2436 33 2450 1122
rect 2464 47 2478 1136
rect 2492 33 2506 1122
rect 2520 47 2534 1136
rect 2548 33 2562 1122
rect 2576 47 2590 1136
rect 2604 33 2618 1122
rect 2632 47 2646 1136
rect 2660 33 2674 1122
rect 2688 47 2702 1136
rect 2716 33 2730 1122
rect 2744 47 2758 1136
rect 2772 33 2786 1122
rect 2800 47 2814 1136
rect 2828 33 2842 1122
rect 2856 47 2870 1136
rect 2884 33 2898 1122
rect 2912 47 2926 1136
rect 2940 33 2954 1122
rect 2968 47 2982 1136
rect 2996 33 3010 1122
rect 3024 47 3038 1136
rect 3052 33 3066 1122
rect 3080 47 3094 1136
rect 3108 33 3122 1122
rect 3136 47 3150 1136
rect 3164 33 3178 1122
rect 3192 47 3206 1136
rect 3220 33 3234 1122
rect 3248 47 3262 1136
rect 3276 33 3290 1122
rect 3304 47 3318 1136
rect 3332 33 3346 1122
rect 3360 47 3374 1136
rect 3388 33 3402 1122
rect 3416 47 3430 1136
rect 3444 33 3458 1122
rect 3472 47 3486 1136
rect 3500 33 3514 1122
rect 3528 47 3542 1136
rect 3556 33 3570 1122
rect 3584 47 3598 1136
rect 3612 33 3626 1122
rect 3640 47 3654 1136
rect 3668 33 3682 1122
rect 3696 47 3710 1136
rect 3724 33 3738 1122
rect 3752 47 3766 1136
rect 3780 33 3794 1122
rect 3808 47 3822 1136
rect 3836 33 3850 1122
rect 3864 47 3878 1136
rect 3892 33 3906 1122
rect 3920 47 3934 1136
rect 3948 33 3962 1122
rect 3976 47 3990 1136
rect 4004 33 4018 1122
rect 4032 47 4046 1136
rect 4060 33 4074 1122
rect 4088 47 4102 1136
rect 4116 33 4130 1122
rect 4144 47 4158 1136
rect 4172 33 4186 1122
rect 4200 47 4214 1136
rect 4228 33 4242 1122
rect 4256 47 4270 1136
rect 4284 33 4298 1122
rect 4312 47 4326 1136
rect 4340 33 4354 1122
rect 4368 47 4382 1136
rect 4396 33 4410 1122
rect 4424 47 4438 1136
rect 4452 33 4466 1122
rect 4480 47 4494 1136
rect 4508 33 4522 1122
rect 4536 47 4550 1136
rect 4564 33 4578 1122
rect 4592 47 4606 1136
rect 4620 33 4634 1122
rect 4648 47 4662 1136
rect 4676 33 4690 1122
rect 4704 47 4718 1136
rect 4732 33 4746 1122
rect 4760 47 4774 1136
rect 4788 33 4802 1122
rect 4816 47 4830 1136
rect 4844 33 4858 1122
rect 4872 47 4886 1136
rect 4900 33 4914 1122
rect 4928 47 4942 1136
rect 4956 33 4970 1122
rect 4984 47 4998 1136
rect 5012 33 5026 1122
rect 5040 47 5054 1136
rect 5068 33 5082 1122
rect 5096 47 5110 1136
rect 5124 33 5138 1122
rect 5152 47 5166 1136
rect 5180 33 5194 1122
rect 5208 47 5222 1136
rect 5236 33 5250 1122
rect 5264 47 5278 1136
rect 5292 33 5306 1122
rect 5320 47 5334 1136
rect 5348 33 5362 1122
rect 5376 47 5390 1136
rect 5404 33 5418 1122
rect 5432 47 5446 1136
rect 5460 33 5474 1122
rect 5488 47 5502 1136
rect 5516 33 5530 1122
rect 5544 47 5573 1136
rect 0 0 5573 33
<< obsm2 >>
rect 0 33 14 1169
rect 28 1136 98 1169
rect 28 47 42 1136
rect 56 33 70 1122
rect 0 0 70 33
rect 84 0 98 1136
rect 112 33 126 1169
rect 140 1136 210 1169
rect 140 47 154 1136
rect 168 33 182 1122
rect 112 0 182 33
rect 196 0 210 1136
rect 224 33 238 1169
rect 252 1136 322 1169
rect 252 47 266 1136
rect 280 33 294 1122
rect 224 0 294 33
rect 308 0 322 1136
rect 336 33 350 1169
rect 364 1136 434 1169
rect 364 47 378 1136
rect 392 33 406 1122
rect 336 0 406 33
rect 420 0 434 1136
rect 448 33 462 1169
rect 476 1136 546 1169
rect 476 47 490 1136
rect 504 33 518 1122
rect 448 0 518 33
rect 532 0 546 1136
rect 560 33 574 1169
rect 588 1136 658 1169
rect 588 47 602 1136
rect 616 33 630 1122
rect 560 0 630 33
rect 644 0 658 1136
rect 672 33 686 1169
rect 700 1136 770 1169
rect 700 47 714 1136
rect 728 33 742 1122
rect 672 0 742 33
rect 756 0 770 1136
rect 784 33 798 1169
rect 812 1136 882 1169
rect 812 47 826 1136
rect 840 33 854 1122
rect 784 0 854 33
rect 868 0 882 1136
rect 896 33 910 1169
rect 924 1136 994 1169
rect 924 47 938 1136
rect 952 33 966 1122
rect 896 0 966 33
rect 980 0 994 1136
rect 1008 33 1022 1169
rect 1036 1136 1106 1169
rect 1036 47 1050 1136
rect 1064 33 1078 1122
rect 1008 0 1078 33
rect 1092 0 1106 1136
rect 1120 33 1134 1169
rect 1148 1136 1218 1169
rect 1148 47 1162 1136
rect 1176 33 1190 1122
rect 1120 0 1190 33
rect 1204 0 1218 1136
rect 1232 33 1246 1169
rect 1260 1136 1330 1169
rect 1260 47 1274 1136
rect 1288 33 1302 1122
rect 1232 0 1302 33
rect 1316 0 1330 1136
rect 1344 33 1358 1169
rect 1372 1136 1442 1169
rect 1372 47 1386 1136
rect 1400 33 1414 1122
rect 1344 0 1414 33
rect 1428 0 1442 1136
rect 1456 33 1470 1169
rect 1484 1136 1554 1169
rect 1484 47 1498 1136
rect 1512 33 1526 1122
rect 1456 0 1526 33
rect 1540 0 1554 1136
rect 1568 33 1582 1169
rect 1596 1136 1666 1169
rect 1596 47 1610 1136
rect 1624 33 1638 1122
rect 1568 0 1638 33
rect 1652 0 1666 1136
rect 1680 33 1694 1169
rect 1708 1136 1778 1169
rect 1708 47 1722 1136
rect 1736 33 1750 1122
rect 1680 0 1750 33
rect 1764 0 1778 1136
rect 1792 33 1806 1169
rect 1820 1136 1890 1169
rect 1820 47 1834 1136
rect 1848 33 1862 1122
rect 1792 0 1862 33
rect 1876 0 1890 1136
rect 1904 33 1918 1169
rect 1932 1136 2002 1169
rect 1932 47 1946 1136
rect 1960 33 1974 1122
rect 1904 0 1974 33
rect 1988 0 2002 1136
rect 2016 33 2030 1169
rect 2044 1136 2114 1169
rect 2044 47 2058 1136
rect 2072 33 2086 1122
rect 2016 0 2086 33
rect 2100 0 2114 1136
rect 2128 33 2142 1169
rect 2156 1136 2226 1169
rect 2156 47 2170 1136
rect 2184 33 2198 1122
rect 2128 0 2198 33
rect 2212 0 2226 1136
rect 2240 33 2254 1169
rect 2268 1136 2338 1169
rect 2268 47 2282 1136
rect 2296 33 2310 1122
rect 2240 0 2310 33
rect 2324 0 2338 1136
rect 2352 33 2366 1169
rect 2380 1136 2450 1169
rect 2380 47 2394 1136
rect 2408 33 2422 1122
rect 2352 0 2422 33
rect 2436 0 2450 1136
rect 2464 33 2478 1169
rect 2492 1136 2562 1169
rect 2492 47 2506 1136
rect 2520 33 2534 1122
rect 2464 0 2534 33
rect 2548 0 2562 1136
rect 2576 33 2590 1169
rect 2604 1136 2674 1169
rect 2604 47 2618 1136
rect 2632 33 2646 1122
rect 2576 0 2646 33
rect 2660 0 2674 1136
rect 2688 33 2702 1169
rect 2716 1136 2786 1169
rect 2716 47 2730 1136
rect 2744 33 2758 1122
rect 2688 0 2758 33
rect 2772 0 2786 1136
rect 2800 33 2814 1169
rect 2828 1136 2898 1169
rect 2828 47 2842 1136
rect 2856 33 2870 1122
rect 2800 0 2870 33
rect 2884 0 2898 1136
rect 2912 33 2926 1169
rect 2940 1136 3010 1169
rect 2940 47 2954 1136
rect 2968 33 2982 1122
rect 2912 0 2982 33
rect 2996 0 3010 1136
rect 3024 33 3038 1169
rect 3052 1136 3122 1169
rect 3052 47 3066 1136
rect 3080 33 3094 1122
rect 3024 0 3094 33
rect 3108 0 3122 1136
rect 3136 33 3150 1169
rect 3164 1136 3234 1169
rect 3164 47 3178 1136
rect 3192 33 3206 1122
rect 3136 0 3206 33
rect 3220 0 3234 1136
rect 3248 33 3262 1169
rect 3276 1136 3346 1169
rect 3276 47 3290 1136
rect 3304 33 3318 1122
rect 3248 0 3318 33
rect 3332 0 3346 1136
rect 3360 33 3374 1169
rect 3388 1136 3458 1169
rect 3388 47 3402 1136
rect 3416 33 3430 1122
rect 3360 0 3430 33
rect 3444 0 3458 1136
rect 3472 33 3486 1169
rect 3500 1136 3570 1169
rect 3500 47 3514 1136
rect 3528 33 3542 1122
rect 3472 0 3542 33
rect 3556 0 3570 1136
rect 3584 33 3598 1169
rect 3612 1136 3682 1169
rect 3612 47 3626 1136
rect 3640 33 3654 1122
rect 3584 0 3654 33
rect 3668 0 3682 1136
rect 3696 33 3710 1169
rect 3724 1136 3794 1169
rect 3724 47 3738 1136
rect 3752 33 3766 1122
rect 3696 0 3766 33
rect 3780 0 3794 1136
rect 3808 33 3822 1169
rect 3836 1136 3906 1169
rect 3836 47 3850 1136
rect 3864 33 3878 1122
rect 3808 0 3878 33
rect 3892 0 3906 1136
rect 3920 33 3934 1169
rect 3948 1136 4018 1169
rect 3948 47 3962 1136
rect 3976 33 3990 1122
rect 3920 0 3990 33
rect 4004 0 4018 1136
rect 4032 33 4046 1169
rect 4060 1136 4130 1169
rect 4060 47 4074 1136
rect 4088 33 4102 1122
rect 4032 0 4102 33
rect 4116 0 4130 1136
rect 4144 33 4158 1169
rect 4172 1136 4242 1169
rect 4172 47 4186 1136
rect 4200 33 4214 1122
rect 4144 0 4214 33
rect 4228 0 4242 1136
rect 4256 33 4270 1169
rect 4284 1136 4354 1169
rect 4284 47 4298 1136
rect 4312 33 4326 1122
rect 4256 0 4326 33
rect 4340 0 4354 1136
rect 4368 33 4382 1169
rect 4396 1136 4466 1169
rect 4396 47 4410 1136
rect 4424 33 4438 1122
rect 4368 0 4438 33
rect 4452 0 4466 1136
rect 4480 33 4494 1169
rect 4508 1136 4578 1169
rect 4508 47 4522 1136
rect 4536 33 4550 1122
rect 4480 0 4550 33
rect 4564 0 4578 1136
rect 4592 33 4606 1169
rect 4620 1136 4690 1169
rect 4620 47 4634 1136
rect 4648 33 4662 1122
rect 4592 0 4662 33
rect 4676 0 4690 1136
rect 4704 33 4718 1169
rect 4732 1136 4802 1169
rect 4732 47 4746 1136
rect 4760 33 4774 1122
rect 4704 0 4774 33
rect 4788 0 4802 1136
rect 4816 33 4830 1169
rect 4844 1136 4914 1169
rect 4844 47 4858 1136
rect 4872 33 4886 1122
rect 4816 0 4886 33
rect 4900 0 4914 1136
rect 4928 33 4942 1169
rect 4956 1136 5026 1169
rect 4956 47 4970 1136
rect 4984 33 4998 1122
rect 4928 0 4998 33
rect 5012 0 5026 1136
rect 5040 33 5054 1169
rect 5068 1136 5138 1169
rect 5068 47 5082 1136
rect 5096 33 5110 1122
rect 5040 0 5110 33
rect 5124 0 5138 1136
rect 5152 33 5166 1169
rect 5180 1136 5250 1169
rect 5180 47 5194 1136
rect 5208 33 5222 1122
rect 5152 0 5222 33
rect 5236 0 5250 1136
rect 5264 33 5278 1169
rect 5292 1136 5362 1169
rect 5292 47 5306 1136
rect 5320 33 5334 1122
rect 5264 0 5334 33
rect 5348 0 5362 1136
rect 5376 33 5390 1169
rect 5404 1136 5573 1169
rect 5404 47 5418 1136
rect 5432 33 5446 1122
rect 5376 0 5446 33
rect 5460 0 5474 1136
rect 5488 33 5502 1122
rect 5516 47 5530 1136
rect 5544 33 5573 1122
rect 5488 0 5573 33
<< obsm3 >>
rect 0 1136 5573 1169
rect 0 63 30 1136
rect 60 33 90 1106
rect 120 63 150 1136
rect 180 33 210 1106
rect 240 63 270 1136
rect 300 33 330 1106
rect 360 63 390 1136
rect 420 33 450 1106
rect 480 63 510 1136
rect 540 33 570 1106
rect 600 63 630 1136
rect 660 33 690 1106
rect 720 63 750 1136
rect 780 33 810 1106
rect 840 63 870 1136
rect 900 33 930 1106
rect 960 63 990 1136
rect 1020 33 1050 1106
rect 1080 63 1110 1136
rect 1140 33 1170 1106
rect 1200 63 1230 1136
rect 1260 33 1290 1106
rect 1320 63 1350 1136
rect 1380 33 1410 1106
rect 1440 63 1470 1136
rect 1500 33 1530 1106
rect 1560 63 1590 1136
rect 1620 33 1650 1106
rect 1680 63 1710 1136
rect 1740 33 1770 1106
rect 1800 63 1830 1136
rect 1860 33 1890 1106
rect 1920 63 1950 1136
rect 1980 33 2010 1106
rect 2040 63 2070 1136
rect 2100 33 2130 1106
rect 2160 63 2190 1136
rect 2220 33 2250 1106
rect 2280 63 2310 1136
rect 2340 33 2370 1106
rect 2400 63 2430 1136
rect 2460 33 2490 1106
rect 2520 63 2550 1136
rect 2580 33 2610 1106
rect 2640 63 2670 1136
rect 2700 33 2730 1106
rect 2760 63 2790 1136
rect 2820 33 2850 1106
rect 2880 63 2910 1136
rect 2940 33 2970 1106
rect 3000 63 3030 1136
rect 3060 33 3090 1106
rect 3120 63 3150 1136
rect 3180 33 3210 1106
rect 3240 63 3270 1136
rect 3300 33 3330 1106
rect 3360 63 3390 1136
rect 3420 33 3450 1106
rect 3480 63 3510 1136
rect 3540 33 3570 1106
rect 3600 63 3630 1136
rect 3660 33 3690 1106
rect 3720 63 3750 1136
rect 3780 33 3810 1106
rect 3840 63 3870 1136
rect 3900 33 3930 1106
rect 3960 63 3990 1136
rect 4020 33 4050 1106
rect 4080 63 4110 1136
rect 4140 33 4170 1106
rect 4200 63 4230 1136
rect 4260 33 4290 1106
rect 4320 63 4350 1136
rect 4380 33 4410 1106
rect 4440 63 4470 1136
rect 4500 33 4530 1106
rect 4560 63 4590 1136
rect 4620 33 4650 1106
rect 4680 63 4710 1136
rect 4740 33 4770 1106
rect 4800 63 4830 1136
rect 4860 33 4890 1106
rect 4920 63 4950 1136
rect 4980 33 5010 1106
rect 5040 63 5070 1136
rect 5100 33 5130 1106
rect 5160 63 5190 1136
rect 5220 33 5250 1106
rect 5280 63 5310 1136
rect 5340 33 5370 1106
rect 5400 63 5430 1136
rect 5460 33 5490 1106
rect 5520 63 5573 1136
rect 0 0 5573 33
<< obsm4 >>
rect 0 1136 5573 1169
rect 0 33 30 1106
rect 60 999 210 1136
rect 60 63 90 999
rect 120 170 150 969
rect 180 200 210 999
rect 240 170 270 1106
rect 120 33 270 170
rect 300 63 330 1136
rect 360 33 390 1106
rect 420 63 450 1136
rect 480 33 510 1106
rect 540 63 570 1136
rect 600 33 630 1106
rect 660 63 690 1136
rect 720 33 750 1106
rect 780 999 930 1136
rect 780 63 810 999
rect 840 170 870 969
rect 900 200 930 999
rect 960 170 990 1106
rect 840 33 990 170
rect 1020 63 1050 1136
rect 1080 33 1110 1106
rect 1140 63 1170 1136
rect 1200 33 1230 1106
rect 1260 63 1290 1136
rect 1320 33 1350 1106
rect 1380 63 1410 1136
rect 1440 33 1470 1106
rect 1500 999 1650 1136
rect 1500 63 1530 999
rect 1560 170 1590 969
rect 1620 200 1650 999
rect 1680 170 1710 1106
rect 1560 33 1710 170
rect 1740 63 1770 1136
rect 1800 33 1830 1106
rect 1860 63 1890 1136
rect 1920 33 1950 1106
rect 1980 63 2010 1136
rect 2040 33 2070 1106
rect 2100 63 2130 1136
rect 2160 33 2190 1106
rect 2220 999 2370 1136
rect 2220 63 2250 999
rect 2280 170 2310 969
rect 2340 200 2370 999
rect 2400 170 2430 1106
rect 2280 33 2430 170
rect 2460 63 2490 1136
rect 2520 33 2550 1106
rect 2580 63 2610 1136
rect 2640 33 2670 1106
rect 2700 63 2730 1136
rect 2760 33 2790 1106
rect 2820 63 2850 1136
rect 2880 33 2910 1106
rect 2940 999 3090 1136
rect 2940 63 2970 999
rect 3000 170 3030 969
rect 3060 200 3090 999
rect 3120 170 3150 1106
rect 3000 33 3150 170
rect 3180 63 3210 1136
rect 3240 33 3270 1106
rect 3300 63 3330 1136
rect 3360 33 3390 1106
rect 3420 63 3450 1136
rect 3480 33 3510 1106
rect 3540 63 3570 1136
rect 3600 33 3630 1106
rect 3660 999 3810 1136
rect 3660 63 3690 999
rect 3720 170 3750 969
rect 3780 200 3810 999
rect 3840 170 3870 1106
rect 3720 33 3870 170
rect 3900 63 3930 1136
rect 3960 33 3990 1106
rect 4020 63 4050 1136
rect 4080 33 4110 1106
rect 4140 63 4170 1136
rect 4200 33 4230 1106
rect 4260 63 4290 1136
rect 4320 33 4350 1106
rect 4380 999 4530 1136
rect 4380 63 4410 999
rect 4440 170 4470 969
rect 4500 200 4530 999
rect 4560 170 4590 1106
rect 4440 33 4590 170
rect 4620 63 4650 1136
rect 4680 33 4710 1106
rect 4740 63 4770 1136
rect 4800 33 4830 1106
rect 4860 63 4890 1136
rect 4920 33 4950 1106
rect 4980 63 5010 1136
rect 5040 33 5070 1106
rect 5100 999 5250 1136
rect 5100 63 5130 999
rect 5160 170 5190 969
rect 5220 200 5250 999
rect 5280 170 5310 1106
rect 5160 33 5310 170
rect 5340 63 5370 1136
rect 5400 33 5430 1106
rect 5460 63 5490 1136
rect 5520 33 5573 1106
rect 0 0 5573 33
<< obsm5 >>
rect 0 969 5493 1129
rect 0 360 160 969
rect 320 200 480 809
rect 640 360 800 969
rect 960 200 1120 809
rect 1280 360 1440 969
rect 1600 200 1760 809
rect 1920 360 2080 969
rect 2240 200 2400 809
rect 2560 360 2720 969
rect 2880 200 3040 809
rect 3200 360 3360 969
rect 3520 200 3680 809
rect 3840 360 4000 969
rect 4160 200 4320 809
rect 4480 360 4640 969
rect 4800 200 4960 809
rect 5120 360 5493 969
rect 0 40 5493 200
<< properties >>
string FIXED_BBOX 0 0 5573 1169
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2155188
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 1999152
<< end >>
