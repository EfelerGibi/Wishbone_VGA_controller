magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< pwell >>
rect 10 76 766 458
<< nmoslvt >>
rect 204 102 254 432
rect 310 102 360 432
rect 416 102 466 432
rect 522 102 572 432
<< ndiff >>
rect 148 420 204 432
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 254 420 310 432
rect 254 386 265 420
rect 299 386 310 420
rect 254 352 310 386
rect 254 318 265 352
rect 299 318 310 352
rect 254 284 310 318
rect 254 250 265 284
rect 299 250 310 284
rect 254 216 310 250
rect 254 182 265 216
rect 299 182 310 216
rect 254 148 310 182
rect 254 114 265 148
rect 299 114 310 148
rect 254 102 310 114
rect 360 420 416 432
rect 360 386 371 420
rect 405 386 416 420
rect 360 352 416 386
rect 360 318 371 352
rect 405 318 416 352
rect 360 284 416 318
rect 360 250 371 284
rect 405 250 416 284
rect 360 216 416 250
rect 360 182 371 216
rect 405 182 416 216
rect 360 148 416 182
rect 360 114 371 148
rect 405 114 416 148
rect 360 102 416 114
rect 466 420 522 432
rect 466 386 477 420
rect 511 386 522 420
rect 466 352 522 386
rect 466 318 477 352
rect 511 318 522 352
rect 466 284 522 318
rect 466 250 477 284
rect 511 250 522 284
rect 466 216 522 250
rect 466 182 477 216
rect 511 182 522 216
rect 466 148 522 182
rect 466 114 477 148
rect 511 114 522 148
rect 466 102 522 114
rect 572 420 628 432
rect 572 386 583 420
rect 617 386 628 420
rect 572 352 628 386
rect 572 318 583 352
rect 617 318 628 352
rect 572 284 628 318
rect 572 250 583 284
rect 617 250 628 284
rect 572 216 628 250
rect 572 182 583 216
rect 617 182 628 216
rect 572 148 628 182
rect 572 114 583 148
rect 617 114 628 148
rect 572 102 628 114
<< ndiffc >>
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 265 386 299 420
rect 265 318 299 352
rect 265 250 299 284
rect 265 182 299 216
rect 265 114 299 148
rect 371 386 405 420
rect 371 318 405 352
rect 371 250 405 284
rect 371 182 405 216
rect 371 114 405 148
rect 477 386 511 420
rect 477 318 511 352
rect 477 250 511 284
rect 477 182 511 216
rect 477 114 511 148
rect 583 386 617 420
rect 583 318 617 352
rect 583 250 617 284
rect 583 182 617 216
rect 583 114 617 148
<< psubdiff >>
rect 36 386 94 432
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 682 386 740 432
rect 682 352 694 386
rect 728 352 740 386
rect 682 318 740 352
rect 682 284 694 318
rect 728 284 740 318
rect 682 250 740 284
rect 682 216 694 250
rect 728 216 740 250
rect 682 182 740 216
rect 682 148 694 182
rect 728 148 740 182
rect 682 102 740 148
<< psubdiffcont >>
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 694 352 728 386
rect 694 284 728 318
rect 694 216 728 250
rect 694 148 728 182
<< poly >>
rect 185 504 591 524
rect 185 470 201 504
rect 235 470 269 504
rect 303 470 337 504
rect 371 470 405 504
rect 439 470 473 504
rect 507 470 541 504
rect 575 470 591 504
rect 185 454 591 470
rect 204 432 254 454
rect 310 432 360 454
rect 416 432 466 454
rect 522 432 572 454
rect 204 80 254 102
rect 310 80 360 102
rect 416 80 466 102
rect 522 80 572 102
rect 185 64 591 80
rect 185 30 201 64
rect 235 30 269 64
rect 303 30 337 64
rect 371 30 405 64
rect 439 30 473 64
rect 507 30 541 64
rect 575 30 591 64
rect 185 10 591 30
<< polycont >>
rect 201 470 235 504
rect 269 470 303 504
rect 337 470 371 504
rect 405 470 439 504
rect 473 470 507 504
rect 541 470 575 504
rect 201 30 235 64
rect 269 30 303 64
rect 337 30 371 64
rect 405 30 439 64
rect 473 30 507 64
rect 541 30 575 64
<< locali >>
rect 185 470 192 504
rect 235 470 264 504
rect 303 470 336 504
rect 371 470 405 504
rect 442 470 473 504
rect 514 470 541 504
rect 586 470 591 504
rect 159 420 193 436
rect 48 392 82 402
rect 48 320 82 352
rect 48 250 82 284
rect 48 182 82 214
rect 48 132 82 142
rect 159 352 193 358
rect 159 284 193 286
rect 159 248 193 250
rect 159 176 193 182
rect 159 98 193 114
rect 265 420 299 436
rect 265 352 299 358
rect 265 284 299 286
rect 265 248 299 250
rect 265 176 299 182
rect 265 98 299 114
rect 371 420 405 436
rect 371 352 405 358
rect 371 284 405 286
rect 371 248 405 250
rect 371 176 405 182
rect 371 98 405 114
rect 477 420 511 436
rect 477 352 511 358
rect 477 284 511 286
rect 477 248 511 250
rect 477 176 511 182
rect 477 98 511 114
rect 583 420 617 436
rect 583 352 617 358
rect 583 284 617 286
rect 583 248 617 250
rect 583 176 617 182
rect 694 392 728 402
rect 694 320 728 352
rect 694 250 728 284
rect 694 182 728 214
rect 694 132 728 142
rect 583 98 617 114
rect 185 30 192 64
rect 235 30 264 64
rect 303 30 336 64
rect 371 30 405 64
rect 442 30 473 64
rect 514 30 541 64
rect 586 30 591 64
<< viali >>
rect 192 470 201 504
rect 201 470 226 504
rect 264 470 269 504
rect 269 470 298 504
rect 336 470 337 504
rect 337 470 370 504
rect 408 470 439 504
rect 439 470 442 504
rect 480 470 507 504
rect 507 470 514 504
rect 552 470 575 504
rect 575 470 586 504
rect 48 386 82 392
rect 48 358 82 386
rect 48 318 82 320
rect 48 286 82 318
rect 48 216 82 248
rect 48 214 82 216
rect 48 148 82 176
rect 48 142 82 148
rect 159 386 193 392
rect 159 358 193 386
rect 159 318 193 320
rect 159 286 193 318
rect 159 216 193 248
rect 159 214 193 216
rect 159 148 193 176
rect 159 142 193 148
rect 265 386 299 392
rect 265 358 299 386
rect 265 318 299 320
rect 265 286 299 318
rect 265 216 299 248
rect 265 214 299 216
rect 265 148 299 176
rect 265 142 299 148
rect 371 386 405 392
rect 371 358 405 386
rect 371 318 405 320
rect 371 286 405 318
rect 371 216 405 248
rect 371 214 405 216
rect 371 148 405 176
rect 371 142 405 148
rect 477 386 511 392
rect 477 358 511 386
rect 477 318 511 320
rect 477 286 511 318
rect 477 216 511 248
rect 477 214 511 216
rect 477 148 511 176
rect 477 142 511 148
rect 583 386 617 392
rect 583 358 617 386
rect 583 318 617 320
rect 583 286 617 318
rect 583 216 617 248
rect 583 214 617 216
rect 583 148 617 176
rect 583 142 617 148
rect 694 386 728 392
rect 694 358 728 386
rect 694 318 728 320
rect 694 286 728 318
rect 694 216 728 248
rect 694 214 728 216
rect 694 148 728 176
rect 694 142 728 148
rect 192 30 201 64
rect 201 30 226 64
rect 264 30 269 64
rect 269 30 298 64
rect 336 30 337 64
rect 337 30 370 64
rect 408 30 439 64
rect 439 30 442 64
rect 480 30 507 64
rect 507 30 514 64
rect 552 30 575 64
rect 575 30 586 64
<< metal1 >>
rect 180 504 598 524
rect 180 470 192 504
rect 226 470 264 504
rect 298 470 336 504
rect 370 470 408 504
rect 442 470 480 504
rect 514 470 552 504
rect 586 470 598 504
rect 180 458 598 470
rect 36 392 94 420
rect 36 358 48 392
rect 82 358 94 392
rect 36 320 94 358
rect 36 286 48 320
rect 82 286 94 320
rect 36 248 94 286
rect 36 214 48 248
rect 82 214 94 248
rect 36 176 94 214
rect 36 142 48 176
rect 82 142 94 176
rect 36 114 94 142
rect 150 392 202 420
rect 150 358 159 392
rect 193 358 202 392
rect 150 320 202 358
rect 150 286 159 320
rect 193 286 202 320
rect 150 248 202 286
rect 150 236 159 248
rect 193 236 202 248
rect 150 176 202 184
rect 150 172 159 176
rect 193 172 202 176
rect 150 114 202 120
rect 256 414 308 420
rect 256 358 265 362
rect 299 358 308 362
rect 256 350 308 358
rect 256 286 265 298
rect 299 286 308 298
rect 256 248 308 286
rect 256 214 265 248
rect 299 214 308 248
rect 256 176 308 214
rect 256 142 265 176
rect 299 142 308 176
rect 256 114 308 142
rect 362 392 414 420
rect 362 358 371 392
rect 405 358 414 392
rect 362 320 414 358
rect 362 286 371 320
rect 405 286 414 320
rect 362 248 414 286
rect 362 236 371 248
rect 405 236 414 248
rect 362 176 414 184
rect 362 172 371 176
rect 405 172 414 176
rect 362 114 414 120
rect 468 414 520 420
rect 468 358 477 362
rect 511 358 520 362
rect 468 350 520 358
rect 468 286 477 298
rect 511 286 520 298
rect 468 248 520 286
rect 468 214 477 248
rect 511 214 520 248
rect 468 176 520 214
rect 468 142 477 176
rect 511 142 520 176
rect 468 114 520 142
rect 574 392 626 420
rect 574 358 583 392
rect 617 358 626 392
rect 574 320 626 358
rect 574 286 583 320
rect 617 286 626 320
rect 574 248 626 286
rect 574 236 583 248
rect 617 236 626 248
rect 574 176 626 184
rect 574 172 583 176
rect 617 172 626 176
rect 574 114 626 120
rect 682 392 740 420
rect 682 358 694 392
rect 728 358 740 392
rect 682 320 740 358
rect 682 286 694 320
rect 728 286 740 320
rect 682 248 740 286
rect 682 214 694 248
rect 728 214 740 248
rect 682 176 740 214
rect 682 142 694 176
rect 728 142 740 176
rect 682 114 740 142
rect 180 64 598 76
rect 180 30 192 64
rect 226 30 264 64
rect 298 30 336 64
rect 370 30 408 64
rect 442 30 480 64
rect 514 30 552 64
rect 586 30 598 64
rect 180 10 598 30
<< via1 >>
rect 150 214 159 236
rect 159 214 193 236
rect 193 214 202 236
rect 150 184 202 214
rect 150 142 159 172
rect 159 142 193 172
rect 193 142 202 172
rect 150 120 202 142
rect 256 392 308 414
rect 256 362 265 392
rect 265 362 299 392
rect 299 362 308 392
rect 256 320 308 350
rect 256 298 265 320
rect 265 298 299 320
rect 299 298 308 320
rect 362 214 371 236
rect 371 214 405 236
rect 405 214 414 236
rect 362 184 414 214
rect 362 142 371 172
rect 371 142 405 172
rect 405 142 414 172
rect 362 120 414 142
rect 468 392 520 414
rect 468 362 477 392
rect 477 362 511 392
rect 511 362 520 392
rect 468 320 520 350
rect 468 298 477 320
rect 477 298 511 320
rect 511 298 520 320
rect 574 214 583 236
rect 583 214 617 236
rect 617 214 626 236
rect 574 184 626 214
rect 574 142 583 172
rect 583 142 617 172
rect 617 142 626 172
rect 574 120 626 142
<< metal2 >>
rect 10 414 766 420
rect 10 362 256 414
rect 308 362 468 414
rect 520 362 766 414
rect 10 350 766 362
rect 10 298 256 350
rect 308 298 468 350
rect 520 298 766 350
rect 10 292 766 298
rect 10 236 766 242
rect 10 184 150 236
rect 202 184 362 236
rect 414 184 574 236
rect 626 184 766 236
rect 10 172 766 184
rect 10 120 150 172
rect 202 120 362 172
rect 414 120 574 172
rect 626 120 766 172
rect 10 114 766 120
<< labels >>
flabel metal2 s 10 292 30 420 7 FreeSans 300 180 0 0 DRAIN
port 2 nsew
flabel metal2 s 10 114 30 242 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal1 s 180 458 598 524 0 FreeSans 300 0 0 0 GATE
port 4 nsew
flabel metal1 s 682 114 740 130 3 FreeSans 300 90 0 0 SUBSTRATE
port 5 nsew
flabel metal1 s 36 114 94 130 3 FreeSans 300 90 0 0 SUBSTRATE
port 5 nsew
flabel metal1 s 180 10 598 76 0 FreeSans 300 0 0 0 GATE
port 4 nsew
<< properties >>
string GDS_END 6036008
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 6025164
<< end >>
