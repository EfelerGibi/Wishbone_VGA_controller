magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1 157 439 203
rect 1538 157 2006 203
rect 1 21 2006 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 431 47 461 131
rect 526 47 556 131
rect 628 47 658 131
rect 712 47 742 131
rect 796 47 826 131
rect 984 47 1014 131
rect 1068 47 1098 131
rect 1152 47 1182 131
rect 1241 47 1271 131
rect 1349 47 1379 131
rect 1421 47 1451 131
rect 1517 47 1547 131
rect 1624 47 1654 177
rect 1724 47 1754 177
rect 1808 47 1838 177
rect 1892 47 1922 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 426 371 456 497
rect 515 371 545 497
rect 628 369 658 497
rect 712 369 742 497
rect 796 369 826 497
rect 984 369 1014 497
rect 1068 369 1098 497
rect 1152 369 1182 497
rect 1241 369 1271 497
rect 1326 369 1356 497
rect 1421 371 1451 497
rect 1529 371 1559 497
rect 1624 297 1654 497
rect 1708 297 1738 497
rect 1808 297 1838 497
rect 1892 297 1922 497
<< ndiff >>
rect 27 97 79 177
rect 27 63 35 97
rect 69 63 79 97
rect 27 47 79 63
rect 109 165 163 177
rect 109 131 119 165
rect 153 131 163 165
rect 109 97 163 131
rect 109 63 119 97
rect 153 63 163 97
rect 109 47 163 63
rect 193 97 247 177
rect 193 63 203 97
rect 237 63 247 97
rect 193 47 247 63
rect 277 97 331 177
rect 277 63 287 97
rect 321 63 331 97
rect 277 47 331 63
rect 361 131 413 177
rect 1564 131 1624 177
rect 361 93 431 131
rect 361 59 387 93
rect 421 59 431 93
rect 361 47 431 59
rect 461 47 526 131
rect 556 106 628 131
rect 556 72 584 106
rect 618 72 628 106
rect 556 47 628 72
rect 658 106 712 131
rect 658 72 668 106
rect 702 72 712 106
rect 658 47 712 72
rect 742 89 796 131
rect 742 55 752 89
rect 786 55 796 89
rect 742 47 796 55
rect 826 106 878 131
rect 826 72 836 106
rect 870 72 878 106
rect 826 47 878 72
rect 932 98 984 131
rect 932 64 940 98
rect 974 64 984 98
rect 932 47 984 64
rect 1014 106 1068 131
rect 1014 72 1024 106
rect 1058 72 1068 106
rect 1014 47 1068 72
rect 1098 89 1152 131
rect 1098 55 1108 89
rect 1142 55 1152 89
rect 1098 47 1152 55
rect 1182 106 1241 131
rect 1182 72 1192 106
rect 1226 72 1241 106
rect 1182 47 1241 72
rect 1271 101 1349 131
rect 1271 67 1293 101
rect 1327 67 1349 101
rect 1271 47 1349 67
rect 1379 47 1421 131
rect 1451 47 1517 131
rect 1547 89 1624 131
rect 1547 55 1557 89
rect 1591 55 1624 89
rect 1547 47 1624 55
rect 1654 165 1724 177
rect 1654 131 1680 165
rect 1714 131 1724 165
rect 1654 97 1724 131
rect 1654 63 1680 97
rect 1714 63 1724 97
rect 1654 47 1724 63
rect 1754 97 1808 177
rect 1754 63 1764 97
rect 1798 63 1808 97
rect 1754 47 1808 63
rect 1838 165 1892 177
rect 1838 131 1848 165
rect 1882 131 1892 165
rect 1838 97 1892 131
rect 1838 63 1848 97
rect 1882 63 1892 97
rect 1838 47 1892 63
rect 1922 97 1980 177
rect 1922 63 1932 97
rect 1966 63 1980 97
rect 1922 47 1980 63
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 297 79 375
rect 109 477 163 497
rect 109 443 119 477
rect 153 443 163 477
rect 109 409 163 443
rect 109 375 119 409
rect 153 375 163 409
rect 109 341 163 375
rect 109 307 119 341
rect 153 307 163 341
rect 109 297 163 307
rect 193 477 247 497
rect 193 443 203 477
rect 237 443 247 477
rect 193 409 247 443
rect 193 375 203 409
rect 237 375 247 409
rect 193 297 247 375
rect 277 477 331 497
rect 277 443 287 477
rect 321 443 331 477
rect 277 409 331 443
rect 277 375 287 409
rect 321 375 331 409
rect 277 297 331 375
rect 361 489 426 497
rect 361 455 379 489
rect 413 455 426 489
rect 361 371 426 455
rect 456 371 515 497
rect 545 484 628 497
rect 545 450 571 484
rect 605 450 628 484
rect 545 416 628 450
rect 545 382 571 416
rect 605 382 628 416
rect 545 371 628 382
rect 361 297 411 371
rect 569 369 628 371
rect 658 456 712 497
rect 658 422 668 456
rect 702 422 712 456
rect 658 369 712 422
rect 742 489 796 497
rect 742 455 752 489
rect 786 455 796 489
rect 742 369 796 455
rect 826 456 878 497
rect 826 422 836 456
rect 870 422 878 456
rect 826 369 878 422
rect 932 485 984 497
rect 932 451 940 485
rect 974 451 984 485
rect 932 417 984 451
rect 932 383 940 417
rect 974 383 984 417
rect 932 369 984 383
rect 1014 472 1068 497
rect 1014 438 1024 472
rect 1058 438 1068 472
rect 1014 369 1068 438
rect 1098 489 1152 497
rect 1098 455 1108 489
rect 1142 455 1152 489
rect 1098 369 1152 455
rect 1182 472 1241 497
rect 1182 438 1192 472
rect 1226 438 1241 472
rect 1182 369 1241 438
rect 1271 477 1326 497
rect 1271 443 1282 477
rect 1316 443 1326 477
rect 1271 369 1326 443
rect 1356 371 1421 497
rect 1451 371 1529 497
rect 1559 489 1624 497
rect 1559 455 1579 489
rect 1613 455 1624 489
rect 1559 371 1624 455
rect 1356 369 1406 371
rect 1574 297 1624 371
rect 1654 477 1708 497
rect 1654 443 1664 477
rect 1698 443 1708 477
rect 1654 409 1708 443
rect 1654 375 1664 409
rect 1698 375 1708 409
rect 1654 297 1708 375
rect 1738 477 1808 497
rect 1738 443 1748 477
rect 1782 443 1808 477
rect 1738 409 1808 443
rect 1738 375 1748 409
rect 1782 375 1808 409
rect 1738 297 1808 375
rect 1838 477 1892 497
rect 1838 443 1848 477
rect 1882 443 1892 477
rect 1838 409 1892 443
rect 1838 375 1848 409
rect 1882 375 1892 409
rect 1838 341 1892 375
rect 1838 307 1848 341
rect 1882 307 1892 341
rect 1838 297 1892 307
rect 1922 477 1981 497
rect 1922 443 1932 477
rect 1966 443 1981 477
rect 1922 409 1981 443
rect 1922 375 1932 409
rect 1966 375 1981 409
rect 1922 297 1981 375
<< ndiffc >>
rect 35 63 69 97
rect 119 131 153 165
rect 119 63 153 97
rect 203 63 237 97
rect 287 63 321 97
rect 387 59 421 93
rect 584 72 618 106
rect 668 72 702 106
rect 752 55 786 89
rect 836 72 870 106
rect 940 64 974 98
rect 1024 72 1058 106
rect 1108 55 1142 89
rect 1192 72 1226 106
rect 1293 67 1327 101
rect 1557 55 1591 89
rect 1680 131 1714 165
rect 1680 63 1714 97
rect 1764 63 1798 97
rect 1848 131 1882 165
rect 1848 63 1882 97
rect 1932 63 1966 97
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 443 153 477
rect 119 375 153 409
rect 119 307 153 341
rect 203 443 237 477
rect 203 375 237 409
rect 287 443 321 477
rect 287 375 321 409
rect 379 455 413 489
rect 571 450 605 484
rect 571 382 605 416
rect 668 422 702 456
rect 752 455 786 489
rect 836 422 870 456
rect 940 451 974 485
rect 940 383 974 417
rect 1024 438 1058 472
rect 1108 455 1142 489
rect 1192 438 1226 472
rect 1282 443 1316 477
rect 1579 455 1613 489
rect 1664 443 1698 477
rect 1664 375 1698 409
rect 1748 443 1782 477
rect 1748 375 1782 409
rect 1848 443 1882 477
rect 1848 375 1882 409
rect 1848 307 1882 341
rect 1932 443 1966 477
rect 1932 375 1966 409
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 426 497 456 523
rect 515 497 545 523
rect 628 497 658 523
rect 712 497 742 523
rect 796 497 826 523
rect 984 497 1014 523
rect 1068 497 1098 523
rect 1152 497 1182 523
rect 1241 497 1271 523
rect 1326 497 1356 523
rect 1421 497 1451 523
rect 1529 497 1559 523
rect 1624 497 1654 523
rect 1708 497 1738 523
rect 1808 497 1838 523
rect 1892 497 1922 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 331 265 361 297
rect 426 265 456 371
rect 515 339 545 371
rect 502 323 556 339
rect 502 289 512 323
rect 546 289 556 323
rect 502 273 556 289
rect 79 249 361 265
rect 79 215 137 249
rect 171 215 205 249
rect 239 215 273 249
rect 307 215 361 249
rect 79 199 361 215
rect 406 249 460 265
rect 406 215 416 249
rect 450 229 460 249
rect 450 215 461 229
rect 406 199 461 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 331 177 361 199
rect 431 131 461 199
rect 526 131 556 273
rect 628 271 658 369
rect 712 272 742 369
rect 796 354 826 369
rect 984 354 1014 369
rect 796 324 1014 354
rect 1068 337 1098 369
rect 939 321 1014 324
rect 939 287 949 321
rect 983 287 1014 321
rect 616 255 670 271
rect 616 221 626 255
rect 660 221 670 255
rect 616 205 670 221
rect 712 256 766 272
rect 939 271 1014 287
rect 1056 321 1110 337
rect 1056 287 1066 321
rect 1100 287 1110 321
rect 1056 271 1110 287
rect 712 222 722 256
rect 756 222 766 256
rect 712 206 766 222
rect 628 131 658 205
rect 712 131 742 206
rect 984 176 1014 271
rect 1069 176 1099 271
rect 1152 241 1182 369
rect 1241 241 1271 369
rect 1326 337 1356 369
rect 1421 339 1451 371
rect 1325 321 1379 337
rect 1325 287 1335 321
rect 1369 287 1379 321
rect 1325 271 1379 287
rect 796 146 1014 176
rect 796 131 826 146
rect 984 131 1014 146
rect 1068 146 1099 176
rect 1141 225 1195 241
rect 1141 191 1151 225
rect 1185 191 1195 225
rect 1141 175 1195 191
rect 1241 225 1295 241
rect 1241 191 1251 225
rect 1285 191 1295 225
rect 1241 175 1295 191
rect 1068 131 1098 146
rect 1152 131 1182 175
rect 1241 131 1271 175
rect 1349 131 1379 271
rect 1421 323 1475 339
rect 1421 289 1431 323
rect 1465 289 1475 323
rect 1421 273 1475 289
rect 1421 131 1451 273
rect 1529 265 1559 371
rect 1624 265 1654 297
rect 1708 265 1738 297
rect 1808 265 1838 297
rect 1892 265 1922 297
rect 1517 249 1571 265
rect 1517 215 1527 249
rect 1561 215 1571 249
rect 1517 199 1571 215
rect 1624 249 1922 265
rect 1624 215 1635 249
rect 1669 215 1703 249
rect 1737 215 1771 249
rect 1805 215 1839 249
rect 1873 215 1922 249
rect 1624 199 1922 215
rect 1517 131 1547 199
rect 1624 177 1654 199
rect 1724 177 1754 199
rect 1808 177 1838 199
rect 1892 177 1922 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 431 21 461 47
rect 526 21 556 47
rect 628 21 658 47
rect 712 21 742 47
rect 796 21 826 47
rect 984 21 1014 47
rect 1068 21 1098 47
rect 1152 21 1182 47
rect 1241 21 1271 47
rect 1349 21 1379 47
rect 1421 21 1451 47
rect 1517 21 1547 47
rect 1624 21 1654 47
rect 1724 21 1754 47
rect 1808 21 1838 47
rect 1892 21 1922 47
<< polycont >>
rect 512 289 546 323
rect 137 215 171 249
rect 205 215 239 249
rect 273 215 307 249
rect 416 215 450 249
rect 949 287 983 321
rect 626 221 660 255
rect 1066 287 1100 321
rect 722 222 756 256
rect 1335 287 1369 321
rect 1151 191 1185 225
rect 1251 191 1285 225
rect 1431 289 1465 323
rect 1527 215 1561 249
rect 1635 215 1669 249
rect 1703 215 1737 249
rect 1771 215 1805 249
rect 1839 215 1873 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 35 477 69 527
rect 35 409 69 443
rect 35 359 69 375
rect 103 477 169 489
rect 103 443 119 477
rect 153 443 169 477
rect 103 409 169 443
rect 103 375 119 409
rect 153 375 169 409
rect 103 341 169 375
rect 203 477 237 527
rect 203 409 237 443
rect 287 477 329 493
rect 321 443 329 477
rect 363 489 429 527
rect 363 455 379 489
rect 413 455 429 489
rect 547 484 634 493
rect 287 409 329 443
rect 547 450 571 484
rect 605 450 634 484
rect 547 416 634 450
rect 203 359 237 375
rect 280 375 287 390
rect 321 375 329 409
rect 103 317 119 341
rect 17 307 119 317
rect 153 317 169 341
rect 280 356 329 375
rect 428 382 571 416
rect 605 382 634 416
rect 668 456 702 493
rect 736 489 802 527
rect 736 455 752 489
rect 786 455 802 489
rect 836 456 883 493
rect 668 421 702 422
rect 870 422 883 456
rect 836 421 883 422
rect 668 387 883 421
rect 924 485 990 527
rect 924 451 940 485
rect 974 451 990 485
rect 924 417 990 451
rect 924 383 940 417
rect 974 383 990 417
rect 1024 472 1058 493
rect 1092 489 1158 527
rect 1092 455 1108 489
rect 1142 455 1158 489
rect 1192 472 1226 493
rect 1024 421 1058 438
rect 1192 421 1226 438
rect 1282 477 1522 493
rect 1316 443 1522 477
rect 1563 489 1629 527
rect 1563 455 1579 489
rect 1613 455 1629 489
rect 1664 477 1698 493
rect 1282 425 1522 443
rect 1024 387 1226 421
rect 1488 421 1522 425
rect 280 317 314 356
rect 428 333 462 382
rect 355 320 462 333
rect 153 307 314 317
rect 17 283 314 307
rect 348 299 462 320
rect 496 323 616 338
rect 348 286 389 299
rect 496 289 512 323
rect 546 289 582 323
rect 650 314 868 348
rect 17 181 87 283
rect 348 249 382 286
rect 121 215 137 249
rect 171 215 205 249
rect 239 215 273 249
rect 307 215 382 249
rect 17 165 305 181
rect 17 147 119 165
rect 103 131 119 147
rect 153 147 305 165
rect 153 131 169 147
rect 35 97 69 113
rect 35 17 69 63
rect 103 97 169 131
rect 103 63 119 97
rect 153 63 169 97
rect 103 51 169 63
rect 203 97 237 113
rect 271 97 305 147
rect 348 165 382 215
rect 416 255 468 265
rect 650 255 684 314
rect 416 249 490 255
rect 450 221 490 249
rect 524 221 536 255
rect 610 221 626 255
rect 660 221 684 255
rect 722 256 800 272
rect 756 255 800 256
rect 756 222 766 255
rect 722 221 766 222
rect 450 215 536 221
rect 416 199 536 215
rect 722 206 800 221
rect 834 250 868 314
rect 916 323 999 349
rect 1319 337 1369 391
rect 1488 387 1621 421
rect 916 321 954 323
rect 916 287 949 321
rect 988 289 999 323
rect 983 287 999 289
rect 1044 321 1369 337
rect 1044 287 1066 321
rect 1100 303 1335 321
rect 1100 287 1116 303
rect 1319 287 1335 303
rect 1415 323 1552 347
rect 1415 289 1431 323
rect 1465 289 1506 323
rect 1540 289 1552 323
rect 1587 328 1621 387
rect 1664 409 1698 443
rect 1748 477 1782 527
rect 1748 409 1782 443
rect 1698 375 1714 393
rect 1664 359 1714 375
rect 1748 359 1782 375
rect 1832 477 1898 485
rect 1832 443 1848 477
rect 1882 443 1898 477
rect 1832 409 1898 443
rect 1832 375 1848 409
rect 1882 375 1898 409
rect 1587 294 1645 328
rect 1044 250 1078 287
rect 1319 271 1369 287
rect 834 193 1078 250
rect 1129 221 1138 255
rect 1172 225 1201 255
rect 1129 191 1151 221
rect 1185 191 1201 225
rect 1235 191 1251 225
rect 1285 191 1372 225
rect 1406 221 1414 255
rect 1448 249 1577 255
rect 1448 221 1527 249
rect 1406 215 1527 221
rect 1561 215 1577 249
rect 1406 199 1577 215
rect 1611 249 1645 294
rect 1680 317 1714 359
rect 1832 341 1898 375
rect 1932 477 1966 527
rect 1932 409 1966 443
rect 1932 359 1966 375
rect 1832 317 1848 341
rect 1680 307 1848 317
rect 1882 317 1898 341
rect 1882 307 2007 317
rect 1680 283 2007 307
rect 1611 215 1635 249
rect 1669 215 1703 249
rect 1737 215 1771 249
rect 1805 215 1839 249
rect 1873 215 1889 249
rect 1269 187 1372 191
rect 570 165 582 187
rect 348 153 582 165
rect 616 153 618 187
rect 348 131 618 153
rect 474 106 618 131
rect 271 63 287 97
rect 321 63 337 97
rect 203 17 237 63
rect 371 59 387 93
rect 421 59 437 93
rect 371 17 437 59
rect 474 72 584 106
rect 474 51 618 72
rect 668 123 870 157
rect 668 106 702 123
rect 836 106 870 123
rect 668 51 702 72
rect 736 55 752 89
rect 786 55 802 89
rect 736 17 802 55
rect 1024 123 1226 157
rect 1269 153 1322 187
rect 1356 153 1372 187
rect 1611 165 1645 215
rect 1940 181 2007 283
rect 1024 106 1058 123
rect 836 51 870 72
rect 924 64 940 98
rect 974 64 990 98
rect 924 17 990 64
rect 1192 106 1226 123
rect 1461 131 1645 165
rect 1680 165 2007 181
rect 1714 147 1848 165
rect 1714 131 1730 147
rect 1024 51 1058 72
rect 1092 55 1108 89
rect 1142 55 1158 89
rect 1092 17 1158 55
rect 1192 51 1226 72
rect 1293 101 1327 119
rect 1461 101 1495 131
rect 1327 67 1495 101
rect 1680 97 1730 131
rect 1832 131 1848 147
rect 1882 147 2007 165
rect 1882 131 1898 147
rect 1293 51 1495 67
rect 1541 55 1557 89
rect 1591 55 1607 89
rect 1541 17 1607 55
rect 1664 63 1680 97
rect 1714 63 1730 97
rect 1664 51 1730 63
rect 1764 97 1798 113
rect 1764 17 1798 63
rect 1832 97 1898 131
rect 1832 63 1848 97
rect 1882 63 1898 97
rect 1832 54 1898 63
rect 1932 97 1966 113
rect 1932 17 1966 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 582 289 616 323
rect 490 221 524 255
rect 766 221 800 255
rect 954 321 988 323
rect 954 289 983 321
rect 983 289 988 321
rect 1506 289 1540 323
rect 1138 225 1172 255
rect 1138 221 1151 225
rect 1151 221 1172 225
rect 1414 221 1448 255
rect 582 153 616 187
rect 1322 153 1356 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 570 323 628 329
rect 570 289 582 323
rect 616 320 628 323
rect 942 323 1000 329
rect 942 320 954 323
rect 616 292 954 320
rect 616 289 628 292
rect 570 283 628 289
rect 942 289 954 292
rect 988 320 1000 323
rect 1494 323 1552 329
rect 1494 320 1506 323
rect 988 292 1506 320
rect 988 289 1000 292
rect 942 283 1000 289
rect 1494 289 1506 292
rect 1540 289 1552 323
rect 1494 283 1552 289
rect 478 255 536 261
rect 478 221 490 255
rect 524 252 536 255
rect 754 255 812 261
rect 754 252 766 255
rect 524 224 766 252
rect 524 221 536 224
rect 478 215 536 221
rect 754 221 766 224
rect 800 252 812 255
rect 1126 255 1184 261
rect 1126 252 1138 255
rect 800 224 1138 252
rect 800 221 812 224
rect 754 215 812 221
rect 1126 221 1138 224
rect 1172 252 1184 255
rect 1402 255 1460 261
rect 1402 252 1414 255
rect 1172 224 1414 252
rect 1172 221 1184 224
rect 1126 215 1184 221
rect 1402 221 1414 224
rect 1448 221 1460 255
rect 1402 215 1460 221
rect 570 187 628 193
rect 570 153 582 187
rect 616 184 628 187
rect 1310 187 1368 193
rect 1310 184 1322 187
rect 616 156 1322 184
rect 616 153 628 156
rect 570 147 628 153
rect 1310 153 1322 156
rect 1356 153 1368 187
rect 1310 147 1368 153
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
flabel locali s 122 357 156 391 0 FreeSans 200 0 0 0 COUT
port 8 nsew signal output
flabel locali s 1966 221 2000 255 0 FreeSans 200 0 0 0 SUM
port 9 nsew signal output
flabel locali s 490 221 524 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 582 289 616 323 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 1322 357 1356 391 0 FreeSans 200 0 0 0 CIN
port 3 nsew signal input
flabel locali s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel locali s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 fa_4
rlabel locali s 722 206 800 272 1 A
port 1 nsew signal input
rlabel locali s 1129 191 1201 255 1 A
port 1 nsew signal input
rlabel locali s 1406 199 1577 255 1 A
port 1 nsew signal input
rlabel metal1 s 1402 252 1460 261 1 A
port 1 nsew signal input
rlabel metal1 s 1402 215 1460 224 1 A
port 1 nsew signal input
rlabel metal1 s 1126 252 1184 261 1 A
port 1 nsew signal input
rlabel metal1 s 1126 215 1184 224 1 A
port 1 nsew signal input
rlabel metal1 s 754 252 812 261 1 A
port 1 nsew signal input
rlabel metal1 s 754 215 812 224 1 A
port 1 nsew signal input
rlabel metal1 s 478 252 536 261 1 A
port 1 nsew signal input
rlabel metal1 s 478 224 1460 252 1 A
port 1 nsew signal input
rlabel metal1 s 478 215 536 224 1 A
port 1 nsew signal input
rlabel locali s 916 287 999 349 1 B
port 2 nsew signal input
rlabel locali s 1415 289 1552 347 1 B
port 2 nsew signal input
rlabel metal1 s 1494 320 1552 329 1 B
port 2 nsew signal input
rlabel metal1 s 1494 283 1552 292 1 B
port 2 nsew signal input
rlabel metal1 s 942 320 1000 329 1 B
port 2 nsew signal input
rlabel metal1 s 942 283 1000 292 1 B
port 2 nsew signal input
rlabel metal1 s 570 320 628 329 1 B
port 2 nsew signal input
rlabel metal1 s 570 292 1552 320 1 B
port 2 nsew signal input
rlabel metal1 s 570 283 628 292 1 B
port 2 nsew signal input
rlabel metal1 s 0 -48 2024 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2024 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2024 544
string GDS_END 2093974
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2078288
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 50.600 0.000 
<< end >>
