magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -66 377 546 897
<< pwell >>
rect 54 43 476 283
rect -26 -43 506 43
<< locali >>
rect 25 355 263 424
rect 299 355 365 424
rect 404 319 455 751
rect 240 285 455 319
rect 240 99 306 285
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 480 831
rect 18 735 352 751
rect 18 701 24 735
rect 58 701 96 735
rect 130 701 168 735
rect 202 701 240 735
rect 274 701 312 735
rect 346 701 352 735
rect 18 460 352 701
rect 18 113 204 265
rect 18 79 22 113
rect 56 79 94 113
rect 128 79 166 113
rect 200 79 204 113
rect 344 113 462 249
rect 18 73 204 79
rect 344 79 350 113
rect 384 79 422 113
rect 456 79 462 113
rect 344 73 462 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 24 701 58 735
rect 96 701 130 735
rect 168 701 202 735
rect 240 701 274 735
rect 312 701 346 735
rect 22 79 56 113
rect 94 79 128 113
rect 166 79 200 113
rect 350 79 384 113
rect 422 79 456 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 831 480 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 480 831
rect 0 791 480 797
rect 0 735 480 763
rect 0 701 24 735
rect 58 701 96 735
rect 130 701 168 735
rect 202 701 240 735
rect 274 701 312 735
rect 346 701 480 735
rect 0 689 480 701
rect 0 113 480 125
rect 0 79 22 113
rect 56 79 94 113
rect 128 79 166 113
rect 200 79 350 113
rect 384 79 422 113
rect 456 79 480 113
rect 0 51 480 79
rect 0 17 480 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -23 480 -17
<< labels >>
rlabel locali s 25 355 263 424 6 A
port 1 nsew signal input
rlabel locali s 299 355 365 424 6 B
port 2 nsew signal input
rlabel metal1 s 0 51 480 125 6 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 -23 480 23 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s -26 -43 506 43 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s 54 43 476 283 6 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 791 480 837 6 VPB
port 5 nsew power bidirectional
rlabel nwell s -66 377 546 897 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 689 480 763 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 240 99 306 285 6 Y
port 7 nsew signal output
rlabel locali s 240 285 455 319 6 Y
port 7 nsew signal output
rlabel locali s 404 319 455 751 6 Y
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 480 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 195320
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 187998
<< end >>
