magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 1 21 911 203
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 167 47 197 177
rect 251 47 281 177
rect 403 47 433 177
rect 511 47 541 177
rect 611 47 641 177
rect 695 47 725 177
rect 803 47 833 177
<< scpmoshvt >>
rect 83 297 113 497
rect 167 297 197 497
rect 251 297 281 497
rect 335 297 365 497
rect 527 297 557 497
rect 611 297 641 497
rect 695 297 725 497
rect 803 297 833 497
<< ndiff >>
rect 27 157 83 177
rect 27 123 39 157
rect 73 123 83 157
rect 27 89 83 123
rect 27 55 39 89
rect 73 55 83 89
rect 27 47 83 55
rect 113 93 167 177
rect 113 59 123 93
rect 157 59 167 93
rect 113 47 167 59
rect 197 157 251 177
rect 197 123 207 157
rect 241 123 251 157
rect 197 89 251 123
rect 197 55 207 89
rect 241 55 251 89
rect 197 47 251 55
rect 281 93 403 177
rect 281 59 291 93
rect 325 59 359 93
rect 393 59 403 93
rect 281 47 403 59
rect 433 157 511 177
rect 433 123 451 157
rect 485 123 511 157
rect 433 89 511 123
rect 433 55 451 89
rect 485 55 511 89
rect 433 47 511 55
rect 541 89 611 177
rect 541 55 551 89
rect 585 55 611 89
rect 541 47 611 55
rect 641 157 695 177
rect 641 123 651 157
rect 685 123 695 157
rect 641 89 695 123
rect 641 55 651 89
rect 685 55 695 89
rect 641 47 695 55
rect 725 168 803 177
rect 725 134 751 168
rect 785 134 803 168
rect 725 47 803 134
rect 833 101 885 177
rect 833 67 843 101
rect 877 67 885 101
rect 833 47 885 67
<< pdiff >>
rect 27 489 83 497
rect 27 455 39 489
rect 73 455 83 489
rect 27 421 83 455
rect 27 387 39 421
rect 73 387 83 421
rect 27 353 83 387
rect 27 319 39 353
rect 73 319 83 353
rect 27 297 83 319
rect 113 485 167 497
rect 113 451 123 485
rect 157 451 167 485
rect 113 417 167 451
rect 113 383 123 417
rect 157 383 167 417
rect 113 297 167 383
rect 197 489 251 497
rect 197 455 207 489
rect 241 455 251 489
rect 197 421 251 455
rect 197 387 207 421
rect 241 387 251 421
rect 197 353 251 387
rect 197 319 207 353
rect 241 319 251 353
rect 197 297 251 319
rect 281 444 335 497
rect 281 410 291 444
rect 325 410 335 444
rect 281 297 335 410
rect 365 421 417 497
rect 365 387 375 421
rect 409 387 417 421
rect 365 353 417 387
rect 365 319 375 353
rect 409 319 417 353
rect 365 297 417 319
rect 471 421 527 497
rect 471 387 483 421
rect 517 387 527 421
rect 471 353 527 387
rect 471 319 483 353
rect 517 319 527 353
rect 471 297 527 319
rect 557 444 611 497
rect 557 410 567 444
rect 601 410 611 444
rect 557 297 611 410
rect 641 489 695 497
rect 641 455 651 489
rect 685 455 695 489
rect 641 421 695 455
rect 641 387 651 421
rect 685 387 695 421
rect 641 353 695 387
rect 641 319 651 353
rect 685 319 695 353
rect 641 297 695 319
rect 725 489 803 497
rect 725 455 751 489
rect 785 455 803 489
rect 725 421 803 455
rect 725 387 751 421
rect 785 387 803 421
rect 725 297 803 387
rect 833 438 885 497
rect 833 404 843 438
rect 877 404 885 438
rect 833 370 885 404
rect 833 336 843 370
rect 877 336 885 370
rect 833 297 885 336
<< ndiffc >>
rect 39 123 73 157
rect 39 55 73 89
rect 123 59 157 93
rect 207 123 241 157
rect 207 55 241 89
rect 291 59 325 93
rect 359 59 393 93
rect 451 123 485 157
rect 451 55 485 89
rect 551 55 585 89
rect 651 123 685 157
rect 651 55 685 89
rect 751 134 785 168
rect 843 67 877 101
<< pdiffc >>
rect 39 455 73 489
rect 39 387 73 421
rect 39 319 73 353
rect 123 451 157 485
rect 123 383 157 417
rect 207 455 241 489
rect 207 387 241 421
rect 207 319 241 353
rect 291 410 325 444
rect 375 387 409 421
rect 375 319 409 353
rect 483 387 517 421
rect 483 319 517 353
rect 567 410 601 444
rect 651 455 685 489
rect 651 387 685 421
rect 651 319 685 353
rect 751 455 785 489
rect 751 387 785 421
rect 843 404 877 438
rect 843 336 877 370
<< poly >>
rect 83 497 113 523
rect 167 497 197 523
rect 251 497 281 523
rect 335 497 365 523
rect 527 497 557 523
rect 611 497 641 523
rect 695 497 725 523
rect 803 497 833 523
rect 83 259 113 297
rect 167 259 197 297
rect 63 249 197 259
rect 63 215 79 249
rect 113 215 147 249
rect 181 215 197 249
rect 63 205 197 215
rect 83 177 113 205
rect 167 177 197 205
rect 251 259 281 297
rect 335 259 365 297
rect 527 259 557 297
rect 611 259 641 297
rect 251 249 433 259
rect 251 215 298 249
rect 332 215 366 249
rect 400 215 433 249
rect 251 205 433 215
rect 507 249 641 259
rect 507 215 523 249
rect 557 215 591 249
rect 625 215 641 249
rect 507 205 641 215
rect 251 177 281 205
rect 403 177 433 205
rect 511 177 541 205
rect 611 177 641 205
rect 695 265 725 297
rect 803 265 833 297
rect 695 249 899 265
rect 695 215 855 249
rect 889 215 899 249
rect 695 199 899 215
rect 695 177 725 199
rect 803 177 833 199
rect 83 21 113 47
rect 167 21 197 47
rect 251 21 281 47
rect 403 21 433 47
rect 511 21 541 47
rect 611 21 641 47
rect 695 21 725 47
rect 803 21 833 47
<< polycont >>
rect 79 215 113 249
rect 147 215 181 249
rect 298 215 332 249
rect 366 215 400 249
rect 523 215 557 249
rect 591 215 625 249
rect 855 215 889 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 18 489 89 493
rect 18 455 39 489
rect 73 455 89 489
rect 18 421 89 455
rect 18 387 39 421
rect 73 387 89 421
rect 18 353 89 387
rect 123 485 157 527
rect 123 417 157 451
rect 123 367 157 383
rect 191 489 257 493
rect 191 455 207 489
rect 241 455 257 489
rect 191 421 257 455
rect 191 387 207 421
rect 241 387 257 421
rect 18 319 39 353
rect 73 333 89 353
rect 191 353 257 387
rect 291 459 601 493
rect 291 444 325 459
rect 567 444 601 459
rect 291 367 325 410
rect 359 421 425 425
rect 359 387 375 421
rect 409 387 425 421
rect 191 333 207 353
rect 73 319 207 333
rect 241 333 257 353
rect 359 353 425 387
rect 359 333 375 353
rect 241 319 375 333
rect 409 319 425 353
rect 18 299 425 319
rect 467 421 533 425
rect 467 387 483 421
rect 517 387 533 421
rect 467 353 533 387
rect 567 367 601 410
rect 635 489 701 493
rect 635 455 651 489
rect 685 455 701 489
rect 635 421 701 455
rect 635 387 651 421
rect 685 387 701 421
rect 467 319 483 353
rect 517 333 533 353
rect 635 353 701 387
rect 735 489 801 527
rect 735 455 751 489
rect 785 455 801 489
rect 735 421 801 455
rect 735 387 751 421
rect 785 387 801 421
rect 735 367 801 387
rect 835 438 903 493
rect 835 404 843 438
rect 877 404 903 438
rect 835 370 903 404
rect 635 333 651 353
rect 517 319 651 333
rect 685 333 701 353
rect 835 336 843 370
rect 877 336 903 370
rect 835 333 903 336
rect 685 319 903 333
rect 467 299 903 319
rect 18 249 248 265
rect 18 215 79 249
rect 113 215 147 249
rect 181 215 248 249
rect 18 211 248 215
rect 282 249 444 265
rect 282 215 298 249
rect 332 215 366 249
rect 400 215 444 249
rect 282 211 444 215
rect 478 249 641 265
rect 478 215 523 249
rect 557 215 591 249
rect 625 215 641 249
rect 478 211 641 215
rect 18 157 701 177
rect 18 123 39 157
rect 73 143 207 157
rect 73 123 89 143
rect 18 89 89 123
rect 191 123 207 143
rect 241 143 451 157
rect 241 123 257 143
rect 18 55 39 89
rect 73 55 89 89
rect 18 51 89 55
rect 123 93 157 109
rect 123 17 157 59
rect 191 89 257 123
rect 435 123 451 143
rect 485 143 651 157
rect 485 123 501 143
rect 191 55 207 89
rect 241 55 257 89
rect 191 51 257 55
rect 291 93 393 109
rect 325 59 359 93
rect 291 17 393 59
rect 435 89 501 123
rect 635 123 651 143
rect 685 123 701 157
rect 435 55 451 89
rect 485 55 501 89
rect 435 51 501 55
rect 535 89 601 109
rect 535 55 551 89
rect 585 55 601 89
rect 535 17 601 55
rect 635 89 701 123
rect 735 168 801 299
rect 735 134 751 168
rect 785 134 801 168
rect 835 249 903 265
rect 835 215 855 249
rect 889 215 903 249
rect 835 151 903 215
rect 735 119 801 134
rect 635 55 651 89
rect 685 85 701 89
rect 835 101 903 117
rect 835 85 843 101
rect 685 67 843 85
rect 877 67 903 101
rect 685 55 903 67
rect 635 51 903 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 858 425 892 459 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 766 289 800 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 766 221 800 255 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 490 357 524 391 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 858 357 892 391 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 766 153 800 187 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 858 153 892 187 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 857 221 891 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 398 221 432 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 o31ai_2
rlabel metal1 s 0 -48 920 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 920 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 1439140
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1430212
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 4.600 0.000 
<< end >>
