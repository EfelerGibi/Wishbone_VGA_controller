magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 1 21 978 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 267 47 297 177
rect 351 47 381 177
rect 435 47 465 177
rect 519 47 549 177
rect 614 47 644 177
rect 698 47 728 177
rect 782 47 812 177
rect 866 47 896 177
<< scpmoshvt >>
rect 79 297 109 497
rect 174 309 204 497
rect 258 309 288 497
rect 342 309 372 497
rect 426 309 456 497
rect 614 297 644 497
rect 698 297 728 497
rect 782 297 812 497
rect 866 297 896 497
<< ndiff >>
rect 27 129 79 177
rect 27 95 35 129
rect 69 95 79 129
rect 27 47 79 95
rect 109 93 161 177
rect 109 59 119 93
rect 153 59 161 93
rect 109 47 161 59
rect 215 129 267 177
rect 215 95 223 129
rect 257 95 267 129
rect 215 47 267 95
rect 297 89 351 177
rect 297 55 307 89
rect 341 55 351 89
rect 297 47 351 55
rect 381 129 435 177
rect 381 95 391 129
rect 425 95 435 129
rect 381 47 435 95
rect 465 89 519 177
rect 465 55 475 89
rect 509 55 519 89
rect 465 47 519 55
rect 549 129 614 177
rect 549 95 565 129
rect 599 95 614 129
rect 549 47 614 95
rect 644 165 698 177
rect 644 131 654 165
rect 688 131 698 165
rect 644 47 698 131
rect 728 90 782 177
rect 728 56 738 90
rect 772 56 782 90
rect 728 47 782 56
rect 812 165 866 177
rect 812 131 822 165
rect 856 131 866 165
rect 812 47 866 131
rect 896 90 952 177
rect 896 56 906 90
rect 940 56 952 90
rect 896 47 952 56
<< pdiff >>
rect 27 448 79 497
rect 27 414 35 448
rect 69 414 79 448
rect 27 380 79 414
rect 27 346 35 380
rect 69 346 79 380
rect 27 297 79 346
rect 109 489 174 497
rect 109 455 119 489
rect 153 455 174 489
rect 109 421 174 455
rect 109 387 119 421
rect 153 387 174 421
rect 109 309 174 387
rect 204 448 258 497
rect 204 414 214 448
rect 248 414 258 448
rect 204 380 258 414
rect 204 346 214 380
rect 248 346 258 380
rect 204 309 258 346
rect 288 489 342 497
rect 288 455 298 489
rect 332 455 342 489
rect 288 421 342 455
rect 288 387 298 421
rect 332 387 342 421
rect 288 309 342 387
rect 372 448 426 497
rect 372 414 382 448
rect 416 414 426 448
rect 372 380 426 414
rect 372 346 382 380
rect 416 346 426 380
rect 372 309 426 346
rect 456 485 508 497
rect 456 451 466 485
rect 500 451 508 485
rect 456 417 508 451
rect 456 383 466 417
rect 500 383 508 417
rect 456 309 508 383
rect 562 448 614 497
rect 562 414 570 448
rect 604 414 614 448
rect 562 380 614 414
rect 562 346 570 380
rect 604 346 614 380
rect 109 297 159 309
rect 562 297 614 346
rect 644 407 698 497
rect 644 373 654 407
rect 688 373 698 407
rect 644 339 698 373
rect 644 305 654 339
rect 688 305 698 339
rect 644 297 698 305
rect 728 448 782 497
rect 728 414 738 448
rect 772 414 782 448
rect 728 380 782 414
rect 728 346 738 380
rect 772 346 782 380
rect 728 297 782 346
rect 812 407 866 497
rect 812 373 822 407
rect 856 373 866 407
rect 812 339 866 373
rect 812 305 822 339
rect 856 305 866 339
rect 812 297 866 305
rect 896 448 948 497
rect 896 414 906 448
rect 940 414 948 448
rect 896 380 948 414
rect 896 346 906 380
rect 940 346 948 380
rect 896 297 948 346
<< ndiffc >>
rect 35 95 69 129
rect 119 59 153 93
rect 223 95 257 129
rect 307 55 341 89
rect 391 95 425 129
rect 475 55 509 89
rect 565 95 599 129
rect 654 131 688 165
rect 738 56 772 90
rect 822 131 856 165
rect 906 56 940 90
<< pdiffc >>
rect 35 414 69 448
rect 35 346 69 380
rect 119 455 153 489
rect 119 387 153 421
rect 214 414 248 448
rect 214 346 248 380
rect 298 455 332 489
rect 298 387 332 421
rect 382 414 416 448
rect 382 346 416 380
rect 466 451 500 485
rect 466 383 500 417
rect 570 414 604 448
rect 570 346 604 380
rect 654 373 688 407
rect 654 305 688 339
rect 738 414 772 448
rect 738 346 772 380
rect 822 373 856 407
rect 822 305 856 339
rect 906 414 940 448
rect 906 346 940 380
<< poly >>
rect 79 497 109 523
rect 174 497 204 523
rect 258 497 288 523
rect 342 497 372 523
rect 426 497 456 523
rect 614 497 644 523
rect 698 497 728 523
rect 782 497 812 523
rect 866 497 896 523
rect 79 265 109 297
rect 174 294 204 309
rect 258 294 288 309
rect 342 294 372 309
rect 426 294 456 309
rect 174 265 456 294
rect 614 265 644 297
rect 698 265 728 297
rect 782 265 812 297
rect 866 265 896 297
rect 22 264 456 265
rect 22 249 204 264
rect 22 215 32 249
rect 66 235 204 249
rect 498 249 552 265
rect 66 215 109 235
rect 498 222 508 249
rect 22 199 109 215
rect 79 177 109 199
rect 267 215 508 222
rect 542 215 552 249
rect 267 199 552 215
rect 614 249 991 265
rect 614 215 947 249
rect 981 215 991 249
rect 614 199 991 215
rect 267 192 549 199
rect 267 177 297 192
rect 351 177 381 192
rect 435 177 465 192
rect 519 177 549 192
rect 614 177 644 199
rect 698 177 728 199
rect 782 177 812 199
rect 866 177 896 199
rect 79 21 109 47
rect 267 21 297 47
rect 351 21 381 47
rect 435 21 465 47
rect 519 21 549 47
rect 614 21 644 47
rect 698 21 728 47
rect 782 21 812 47
rect 866 21 896 47
<< polycont >>
rect 32 215 66 249
rect 508 215 542 249
rect 947 215 981 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 17 448 69 493
rect 17 414 35 448
rect 17 380 69 414
rect 17 346 35 380
rect 103 489 169 527
rect 103 455 119 489
rect 153 455 169 489
rect 103 421 169 455
rect 103 387 119 421
rect 153 387 169 421
rect 103 367 169 387
rect 203 448 248 493
rect 203 414 214 448
rect 203 380 248 414
rect 17 333 69 346
rect 203 346 214 380
rect 282 489 348 527
rect 282 455 298 489
rect 332 455 348 489
rect 282 421 348 455
rect 282 387 298 421
rect 332 387 348 421
rect 282 367 348 387
rect 382 448 416 493
rect 382 380 416 414
rect 203 333 248 346
rect 450 485 528 527
rect 450 451 466 485
rect 500 451 528 485
rect 450 417 528 451
rect 450 383 466 417
rect 500 383 528 417
rect 450 367 528 383
rect 562 459 995 493
rect 562 448 604 459
rect 562 414 570 448
rect 738 448 772 459
rect 562 380 604 414
rect 382 333 416 346
rect 562 346 570 380
rect 562 333 604 346
rect 17 299 169 333
rect 203 299 604 333
rect 638 407 704 415
rect 638 373 654 407
rect 688 373 704 407
rect 638 339 704 373
rect 638 305 654 339
rect 688 305 704 339
rect 906 448 995 459
rect 738 380 772 414
rect 738 330 772 346
rect 806 407 872 415
rect 806 373 822 407
rect 856 373 872 407
rect 806 339 872 373
rect 103 265 169 299
rect 638 296 704 305
rect 806 305 822 339
rect 856 305 872 339
rect 940 414 995 448
rect 906 380 995 414
rect 940 346 995 380
rect 906 330 995 346
rect 806 296 872 305
rect 17 249 69 265
rect 17 215 32 249
rect 66 215 69 249
rect 17 199 69 215
rect 103 249 604 265
rect 103 215 508 249
rect 542 215 604 249
rect 103 199 604 215
rect 103 165 169 199
rect 638 165 872 296
rect 17 131 169 165
rect 203 131 599 165
rect 17 129 69 131
rect 17 95 35 129
rect 203 129 257 131
rect 17 51 69 95
rect 103 93 169 97
rect 103 59 119 93
rect 153 59 169 93
rect 103 17 169 59
rect 203 95 223 129
rect 391 129 425 131
rect 203 51 257 95
rect 291 89 357 97
rect 291 55 307 89
rect 341 55 357 89
rect 291 17 357 55
rect 565 129 599 131
rect 391 51 425 95
rect 459 89 525 97
rect 459 55 475 89
rect 509 55 525 89
rect 459 17 525 55
rect 638 131 654 165
rect 688 131 822 165
rect 856 131 872 165
rect 638 124 872 131
rect 906 249 995 265
rect 906 215 947 249
rect 981 215 995 249
rect 906 124 995 215
rect 565 90 599 95
rect 565 56 738 90
rect 772 56 906 90
rect 940 56 995 90
rect 565 51 995 56
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 766 153 800 187 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 766 221 800 255 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 674 221 708 255 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 674 153 708 187 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 949 153 983 187 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 949 221 983 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 einvn_4
rlabel metal1 s 0 -48 1012 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1012 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_END 2979906
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2972128
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 25.300 13.600 
<< end >>
