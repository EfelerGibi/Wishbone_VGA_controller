* NGSPICE file created from sky130_fd_pr__rf_npn_11v0_W1p00L1p00.ext - technology: sky130A

.subckt sky130_fd_pr__rf_npn_11v0_W1p00L1p00 E B C
X0 C B a_512_512# VSUBS sky130_fd_pr__npn_11v0 area=80.1
**devattr s=37813,302
.ends

