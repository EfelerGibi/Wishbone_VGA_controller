magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 545 163 735 203
rect 1 27 735 163
rect 30 -17 64 27
rect 545 21 735 27
<< locali >>
rect 122 425 532 483
rect 17 151 85 265
rect 304 199 452 323
rect 664 299 719 493
rect 486 199 562 265
rect 685 152 719 299
rect 664 83 719 152
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 312 85 527
rect 119 265 167 384
rect 206 357 532 391
rect 566 367 622 527
rect 206 299 270 357
rect 498 333 532 357
rect 119 199 250 265
rect 498 299 630 333
rect 596 265 630 299
rect 596 199 651 265
rect 17 17 85 117
rect 119 61 168 199
rect 596 165 630 199
rect 313 131 630 165
rect 207 17 273 117
rect 313 61 347 131
rect 382 17 448 97
rect 482 61 516 131
rect 550 17 626 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 486 199 562 265 6 A
port 1 nsew signal input
rlabel locali s 122 425 532 483 6 B
port 2 nsew signal input
rlabel locali s 304 199 452 323 6 C
port 3 nsew signal input
rlabel locali s 17 151 85 265 6 D_N
port 4 nsew signal input
rlabel metal1 s 0 -48 736 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 545 21 735 27 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 30 -17 64 27 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 27 735 163 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 545 163 735 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 664 83 719 152 6 X
port 9 nsew signal output
rlabel locali s 685 152 719 299 6 X
port 9 nsew signal output
rlabel locali s 664 299 719 493 6 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 736 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1075482
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1068258
<< end >>
