magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 1 21 1143 203
rect 30 -17 64 21
<< scnmos >>
rect 80 47 110 177
rect 166 47 196 177
rect 252 47 282 177
rect 338 47 368 177
rect 432 47 462 177
rect 518 47 548 177
rect 604 47 634 177
rect 690 47 720 177
rect 776 47 806 177
rect 862 47 892 177
rect 948 47 978 177
rect 1034 47 1064 177
<< scpmoshvt >>
rect 80 297 110 497
rect 166 297 196 497
rect 252 297 282 497
rect 338 297 368 497
rect 430 297 460 497
rect 518 297 548 497
rect 604 297 634 497
rect 690 297 720 497
rect 776 297 806 497
rect 862 297 892 497
rect 948 297 978 497
rect 1034 297 1064 497
<< ndiff >>
rect 27 161 80 177
rect 27 127 35 161
rect 69 127 80 161
rect 27 93 80 127
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 124 166 177
rect 110 90 121 124
rect 155 90 166 124
rect 110 47 166 90
rect 196 89 252 177
rect 196 55 207 89
rect 241 55 252 89
rect 196 47 252 55
rect 282 169 338 177
rect 282 135 293 169
rect 327 135 338 169
rect 282 101 338 135
rect 282 67 293 101
rect 327 67 338 101
rect 282 47 338 67
rect 368 89 432 177
rect 368 55 387 89
rect 421 55 432 89
rect 368 47 432 55
rect 462 101 518 177
rect 462 67 473 101
rect 507 67 518 101
rect 462 47 518 67
rect 548 169 604 177
rect 548 135 559 169
rect 593 135 604 169
rect 548 47 604 135
rect 634 101 690 177
rect 634 67 645 101
rect 679 67 690 101
rect 634 47 690 67
rect 720 169 776 177
rect 720 135 731 169
rect 765 135 776 169
rect 720 47 776 135
rect 806 157 862 177
rect 806 123 817 157
rect 851 123 862 157
rect 806 89 862 123
rect 806 55 817 89
rect 851 55 862 89
rect 806 47 862 55
rect 892 97 948 177
rect 892 63 903 97
rect 937 63 948 97
rect 892 47 948 63
rect 978 164 1034 177
rect 978 130 989 164
rect 1023 130 1034 164
rect 978 96 1034 130
rect 978 62 989 96
rect 1023 62 1034 96
rect 978 47 1034 62
rect 1064 161 1117 177
rect 1064 127 1075 161
rect 1109 127 1117 161
rect 1064 93 1117 127
rect 1064 59 1075 93
rect 1109 59 1117 93
rect 1064 47 1117 59
<< pdiff >>
rect 28 477 80 497
rect 28 443 36 477
rect 70 443 80 477
rect 28 409 80 443
rect 28 375 36 409
rect 70 375 80 409
rect 28 297 80 375
rect 110 387 166 497
rect 110 353 121 387
rect 155 353 166 387
rect 110 297 166 353
rect 196 489 252 497
rect 196 455 207 489
rect 241 455 252 489
rect 196 297 252 455
rect 282 395 338 497
rect 282 361 293 395
rect 327 361 338 395
rect 282 297 338 361
rect 368 477 430 497
rect 368 443 385 477
rect 419 443 430 477
rect 368 297 430 443
rect 460 489 518 497
rect 460 455 473 489
rect 507 455 518 489
rect 460 297 518 455
rect 548 477 604 497
rect 548 443 559 477
rect 593 443 604 477
rect 548 409 604 443
rect 548 375 559 409
rect 593 375 604 409
rect 548 297 604 375
rect 634 489 690 497
rect 634 455 645 489
rect 679 455 690 489
rect 634 297 690 455
rect 720 477 776 497
rect 720 443 731 477
rect 765 443 776 477
rect 720 409 776 443
rect 720 375 731 409
rect 765 375 776 409
rect 720 297 776 375
rect 806 489 862 497
rect 806 455 817 489
rect 851 455 862 489
rect 806 297 862 455
rect 892 477 948 497
rect 892 443 903 477
rect 937 443 948 477
rect 892 297 948 443
rect 978 489 1034 497
rect 978 455 989 489
rect 1023 455 1034 489
rect 978 297 1034 455
rect 1064 477 1117 497
rect 1064 443 1075 477
rect 1109 443 1117 477
rect 1064 409 1117 443
rect 1064 375 1075 409
rect 1109 375 1117 409
rect 1064 297 1117 375
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 121 90 155 124
rect 207 55 241 89
rect 293 135 327 169
rect 293 67 327 101
rect 387 55 421 89
rect 473 67 507 101
rect 559 135 593 169
rect 645 67 679 101
rect 731 135 765 169
rect 817 123 851 157
rect 817 55 851 89
rect 903 63 937 97
rect 989 130 1023 164
rect 989 62 1023 96
rect 1075 127 1109 161
rect 1075 59 1109 93
<< pdiffc >>
rect 36 443 70 477
rect 36 375 70 409
rect 121 353 155 387
rect 207 455 241 489
rect 293 361 327 395
rect 385 443 419 477
rect 473 455 507 489
rect 559 443 593 477
rect 559 375 593 409
rect 645 455 679 489
rect 731 443 765 477
rect 731 375 765 409
rect 817 455 851 489
rect 903 443 937 477
rect 989 455 1023 489
rect 1075 443 1109 477
rect 1075 375 1109 409
<< poly >>
rect 80 497 110 523
rect 166 497 196 523
rect 252 497 282 523
rect 338 497 368 523
rect 430 497 460 523
rect 518 497 548 523
rect 604 497 634 523
rect 690 497 720 523
rect 776 497 806 523
rect 862 497 892 523
rect 948 497 978 523
rect 1034 497 1064 523
rect 80 265 110 297
rect 166 265 196 297
rect 252 265 282 297
rect 338 265 368 297
rect 430 265 460 297
rect 22 249 368 265
rect 22 215 32 249
rect 66 215 100 249
rect 134 215 168 249
rect 202 215 236 249
rect 270 215 368 249
rect 22 199 368 215
rect 410 249 476 265
rect 410 215 426 249
rect 460 215 476 249
rect 410 199 476 215
rect 518 259 548 297
rect 604 259 634 297
rect 690 259 720 297
rect 776 259 806 297
rect 518 249 806 259
rect 518 215 542 249
rect 576 215 610 249
rect 644 215 678 249
rect 712 215 746 249
rect 780 215 806 249
rect 80 177 110 199
rect 166 177 196 199
rect 252 177 282 199
rect 338 177 368 199
rect 432 177 462 199
rect 518 198 806 215
rect 518 177 548 198
rect 604 177 634 198
rect 690 177 720 198
rect 776 177 806 198
rect 862 265 892 297
rect 948 265 978 297
rect 1034 265 1064 297
rect 862 249 1088 265
rect 862 215 908 249
rect 942 215 976 249
rect 1010 215 1044 249
rect 1078 215 1088 249
rect 862 199 1088 215
rect 862 177 892 199
rect 948 177 978 199
rect 1034 177 1064 199
rect 80 21 110 47
rect 166 21 196 47
rect 252 21 282 47
rect 338 21 368 47
rect 432 21 462 47
rect 518 21 548 47
rect 604 21 634 47
rect 690 21 720 47
rect 776 21 806 47
rect 862 21 892 47
rect 948 21 978 47
rect 1034 21 1064 47
<< polycont >>
rect 32 215 66 249
rect 100 215 134 249
rect 168 215 202 249
rect 236 215 270 249
rect 426 215 460 249
rect 542 215 576 249
rect 610 215 644 249
rect 678 215 712 249
rect 746 215 780 249
rect 908 215 942 249
rect 976 215 1010 249
rect 1044 215 1078 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 36 489 423 493
rect 36 477 207 489
rect 70 455 207 477
rect 241 477 423 489
rect 241 455 385 477
rect 70 443 385 455
rect 419 443 423 477
rect 457 489 523 527
rect 457 455 473 489
rect 507 455 523 489
rect 557 477 595 493
rect 36 409 75 443
rect 191 441 423 443
rect 70 375 75 409
rect 383 421 423 441
rect 557 443 559 477
rect 593 443 595 477
rect 629 489 695 527
rect 629 455 645 489
rect 679 455 695 489
rect 729 477 767 493
rect 557 421 595 443
rect 729 443 731 477
rect 765 443 767 477
rect 801 489 867 527
rect 801 455 817 489
rect 851 455 867 489
rect 901 477 937 493
rect 729 421 767 443
rect 901 443 903 477
rect 973 489 1039 527
rect 973 455 989 489
rect 1023 455 1039 489
rect 1073 477 1125 493
rect 901 421 937 443
rect 1073 443 1075 477
rect 1109 443 1125 477
rect 1073 421 1125 443
rect 383 409 1125 421
rect 36 359 75 375
rect 116 395 349 407
rect 116 387 293 395
rect 116 353 121 387
rect 155 361 293 387
rect 327 361 349 395
rect 383 375 559 409
rect 593 375 731 409
rect 765 375 1075 409
rect 1109 375 1125 409
rect 155 353 349 361
rect 116 341 349 353
rect 116 317 376 341
rect 18 249 286 283
rect 18 215 32 249
rect 66 215 100 249
rect 134 215 168 249
rect 202 215 236 249
rect 270 215 286 249
rect 18 207 286 215
rect 18 199 80 207
rect 320 179 376 317
rect 410 296 1094 341
rect 410 249 479 296
rect 410 215 426 249
rect 460 215 479 249
rect 410 213 479 215
rect 513 249 800 262
rect 513 215 542 249
rect 576 215 610 249
rect 644 215 678 249
rect 712 215 746 249
rect 780 215 800 249
rect 845 249 1094 296
rect 845 215 908 249
rect 942 215 976 249
rect 1010 215 1044 249
rect 1078 215 1094 249
rect 513 213 800 215
rect 320 173 781 179
rect 119 169 781 173
rect 18 127 35 161
rect 69 127 85 161
rect 18 93 85 127
rect 18 59 35 93
rect 69 59 85 93
rect 119 135 293 169
rect 327 139 559 169
rect 327 135 329 139
rect 455 135 559 139
rect 593 135 731 169
rect 765 135 781 169
rect 815 164 1039 181
rect 815 157 989 164
rect 119 124 329 135
rect 119 90 121 124
rect 155 123 329 124
rect 155 90 157 123
rect 119 74 157 90
rect 291 101 329 123
rect 815 123 817 157
rect 851 147 989 157
rect 851 123 867 147
rect 18 17 85 59
rect 191 55 207 89
rect 241 55 257 89
rect 191 17 257 55
rect 291 67 293 101
rect 327 67 329 101
rect 291 51 329 67
rect 367 89 423 105
rect 815 101 867 123
rect 973 130 989 147
rect 1023 130 1039 164
rect 367 55 387 89
rect 421 55 423 89
rect 367 17 423 55
rect 457 67 473 101
rect 507 67 645 101
rect 679 89 867 101
rect 679 67 817 89
rect 457 55 817 67
rect 851 55 867 89
rect 457 51 867 55
rect 901 97 939 113
rect 901 63 903 97
rect 937 63 939 97
rect 901 17 939 63
rect 973 96 1039 130
rect 973 62 989 96
rect 1023 62 1039 96
rect 973 51 1039 62
rect 1073 161 1125 177
rect 1073 127 1075 161
rect 1109 127 1125 161
rect 1073 93 1125 127
rect 1073 59 1075 93
rect 1109 59 1125 93
rect 1073 17 1125 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 214 221 248 255 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 1042 289 1076 323 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 766 221 800 255 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 306 357 340 391 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 a21oi_4
rlabel metal1 s 0 -48 1196 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1196 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_END 4074444
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4065910
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 29.900 0.000 
<< end >>
