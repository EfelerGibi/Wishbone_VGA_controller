magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect 0 168 168 1076
rect 1206 168 1374 1076
rect 0 0 1374 168
<< pwell >>
rect 228 228 1146 802
<< mvnmos >>
rect 412 415 1012 615
<< mvndiff >>
rect 412 660 1012 668
rect 412 626 490 660
rect 524 626 558 660
rect 592 626 626 660
rect 660 626 694 660
rect 728 626 762 660
rect 796 626 830 660
rect 864 626 898 660
rect 932 626 966 660
rect 1000 626 1012 660
rect 412 615 1012 626
rect 412 404 1012 415
rect 412 370 490 404
rect 524 370 558 404
rect 592 370 626 404
rect 660 370 694 404
rect 728 370 762 404
rect 796 370 830 404
rect 864 370 898 404
rect 932 370 966 404
rect 1000 370 1012 404
rect 412 362 1012 370
<< mvndiffc >>
rect 490 626 524 660
rect 558 626 592 660
rect 626 626 660 660
rect 694 626 728 660
rect 762 626 796 660
rect 830 626 864 660
rect 898 626 932 660
rect 966 626 1000 660
rect 490 370 524 404
rect 558 370 592 404
rect 626 370 660 404
rect 694 370 728 404
rect 762 370 796 404
rect 830 370 864 404
rect 898 370 932 404
rect 966 370 1000 404
<< mvpsubdiff >>
rect 254 742 356 776
rect 390 742 424 776
rect 458 742 492 776
rect 526 742 560 776
rect 594 742 628 776
rect 662 742 696 776
rect 730 742 764 776
rect 798 742 832 776
rect 866 742 900 776
rect 934 742 1052 776
rect 254 674 288 708
rect 254 606 288 640
rect 1086 662 1120 776
rect 254 538 288 572
rect 254 470 288 504
rect 254 402 288 436
rect 1086 594 1120 628
rect 1086 526 1120 560
rect 1086 458 1120 492
rect 254 254 288 368
rect 1086 390 1120 424
rect 1086 322 1120 356
rect 322 254 356 288
rect 390 254 424 288
rect 458 254 492 288
rect 526 254 560 288
rect 594 254 628 288
rect 662 254 696 288
rect 730 254 764 288
rect 798 254 832 288
rect 866 254 900 288
rect 934 254 968 288
rect 1002 254 1120 288
<< mvnsubdiff >>
rect 66 909 100 933
rect 66 838 100 875
rect 66 767 100 804
rect 1272 909 1306 933
rect 1272 838 1306 875
rect 66 696 100 733
rect 66 625 100 662
rect 66 554 100 591
rect 66 483 100 520
rect 66 412 100 449
rect 66 341 100 378
rect 66 270 100 307
rect 1272 767 1306 804
rect 1272 696 1306 733
rect 1272 625 1306 662
rect 1272 554 1306 591
rect 1272 483 1306 520
rect 1272 412 1306 449
rect 1272 341 1306 378
rect 1272 270 1306 307
rect 66 199 100 236
rect 66 102 100 165
rect 1272 198 1306 236
rect 1272 126 1306 164
rect 66 68 90 102
rect 124 68 159 102
rect 193 68 228 102
rect 262 68 296 102
rect 330 68 364 102
rect 398 68 432 102
rect 466 68 500 102
rect 534 68 568 102
rect 602 68 636 102
rect 670 68 704 102
rect 738 68 772 102
rect 806 68 840 102
rect 874 68 908 102
rect 942 68 976 102
rect 1010 68 1044 102
rect 1078 68 1112 102
rect 1146 68 1180 102
rect 1214 92 1272 102
rect 1214 68 1306 92
<< mvpsubdiffcont >>
rect 356 742 390 776
rect 424 742 458 776
rect 492 742 526 776
rect 560 742 594 776
rect 628 742 662 776
rect 696 742 730 776
rect 764 742 798 776
rect 832 742 866 776
rect 900 742 934 776
rect 1052 742 1086 776
rect 254 708 288 742
rect 254 640 288 674
rect 1086 628 1120 662
rect 254 572 288 606
rect 254 504 288 538
rect 254 436 288 470
rect 1086 560 1120 594
rect 1086 492 1120 526
rect 1086 424 1120 458
rect 254 368 288 402
rect 1086 356 1120 390
rect 1086 288 1120 322
rect 288 254 322 288
rect 356 254 390 288
rect 424 254 458 288
rect 492 254 526 288
rect 560 254 594 288
rect 628 254 662 288
rect 696 254 730 288
rect 764 254 798 288
rect 832 254 866 288
rect 900 254 934 288
rect 968 254 1002 288
<< mvnsubdiffcont >>
rect 66 875 100 909
rect 66 804 100 838
rect 1272 875 1306 909
rect 1272 804 1306 838
rect 66 733 100 767
rect 66 662 100 696
rect 66 591 100 625
rect 66 520 100 554
rect 66 449 100 483
rect 66 378 100 412
rect 66 307 100 341
rect 66 236 100 270
rect 1272 733 1306 767
rect 1272 662 1306 696
rect 1272 591 1306 625
rect 1272 520 1306 554
rect 1272 449 1306 483
rect 1272 378 1306 412
rect 1272 307 1306 341
rect 66 165 100 199
rect 1272 236 1306 270
rect 1272 164 1306 198
rect 90 68 124 102
rect 159 68 193 102
rect 228 68 262 102
rect 296 68 330 102
rect 364 68 398 102
rect 432 68 466 102
rect 500 68 534 102
rect 568 68 602 102
rect 636 68 670 102
rect 704 68 738 102
rect 772 68 806 102
rect 840 68 874 102
rect 908 68 942 102
rect 976 68 1010 102
rect 1044 68 1078 102
rect 1112 68 1146 102
rect 1180 68 1214 102
rect 1272 92 1306 126
<< poly >>
rect 320 599 412 615
rect 320 565 336 599
rect 370 565 412 599
rect 320 531 412 565
rect 320 497 336 531
rect 370 497 412 531
rect 320 463 412 497
rect 320 429 336 463
rect 370 429 412 463
rect 320 415 412 429
rect 1012 415 1038 615
rect 320 413 386 415
<< polycont >>
rect 336 565 370 599
rect 336 497 370 531
rect 336 429 370 463
<< locali >>
rect 877 5301 915 5335
rect 949 5301 987 5335
rect 66 909 100 933
rect 1272 909 1306 933
rect 66 844 68 875
rect 66 838 102 844
rect 100 806 102 838
rect 66 772 68 804
rect 1272 838 1306 841
rect 1272 803 1306 804
rect 66 767 102 772
rect 100 734 102 767
rect 66 700 68 733
rect 66 696 102 700
rect 100 662 102 696
rect 66 628 68 662
rect 66 625 102 628
rect 100 591 102 625
rect 66 590 102 591
rect 66 556 68 590
rect 66 554 102 556
rect 100 520 102 554
rect 66 518 102 520
rect 66 484 68 518
rect 66 483 102 484
rect 100 449 102 483
rect 66 446 102 449
rect 66 412 68 446
rect 100 378 102 412
rect 66 374 102 378
rect 66 341 68 374
rect 100 307 102 340
rect 66 302 102 307
rect 66 270 68 302
rect 100 236 102 268
rect 254 742 276 776
rect 310 742 348 776
rect 390 742 420 776
rect 458 742 492 776
rect 526 742 560 776
rect 598 742 628 776
rect 670 742 696 776
rect 742 742 764 776
rect 814 742 832 776
rect 886 742 900 776
rect 958 742 996 776
rect 1030 742 1052 776
rect 1102 742 1120 776
rect 254 686 288 708
rect 1086 681 1120 742
rect 254 606 288 640
rect 474 626 475 660
rect 524 626 547 660
rect 592 626 619 660
rect 660 626 691 660
rect 728 626 762 660
rect 797 626 830 660
rect 869 626 898 660
rect 941 626 966 660
rect 1013 626 1016 660
rect 254 538 288 570
rect 254 470 288 488
rect 336 599 370 615
rect 336 531 370 538
rect 336 463 370 466
rect 336 413 370 429
rect 1086 609 1120 628
rect 1086 537 1120 560
rect 1086 465 1120 492
rect 254 402 288 407
rect 524 370 556 404
rect 592 370 626 404
rect 671 370 694 404
rect 752 370 762 404
rect 796 370 799 404
rect 864 370 880 404
rect 932 370 961 404
rect 1000 370 1016 404
rect 1086 393 1120 424
rect 254 360 288 368
rect 254 254 288 326
rect 1086 322 1120 356
rect 334 254 356 288
rect 413 254 424 288
rect 526 254 537 288
rect 594 254 616 288
rect 662 254 695 288
rect 730 254 764 288
rect 808 254 832 288
rect 886 254 900 288
rect 964 254 968 288
rect 1002 254 1008 288
rect 1042 254 1086 288
rect 1272 767 1306 769
rect 1272 731 1306 733
rect 1272 696 1306 697
rect 1272 659 1306 662
rect 1272 587 1306 591
rect 1272 515 1306 520
rect 1272 443 1306 449
rect 1272 371 1306 378
rect 1272 299 1306 307
rect 66 230 102 236
rect 66 199 68 230
rect 100 165 102 196
rect 66 158 102 165
rect 66 124 68 158
rect 66 102 102 124
rect 1272 227 1306 236
rect 1272 155 1306 164
rect 66 68 90 102
rect 124 68 138 102
rect 193 68 212 102
rect 262 68 286 102
rect 330 68 360 102
rect 398 68 432 102
rect 468 68 500 102
rect 542 68 568 102
rect 616 68 636 102
rect 690 68 704 102
rect 764 68 772 102
rect 838 68 840 102
rect 874 68 878 102
rect 942 68 952 102
rect 1010 68 1026 102
rect 1078 68 1100 102
rect 1146 68 1174 102
rect 1214 92 1272 102
rect 1214 68 1306 92
<< viali >>
rect 843 5301 877 5335
rect 915 5301 949 5335
rect 987 5301 1021 5335
rect 68 875 100 878
rect 100 875 102 878
rect 68 844 102 875
rect 68 804 100 806
rect 100 804 102 806
rect 68 772 102 804
rect 1272 841 1306 875
rect 68 733 100 734
rect 100 733 102 734
rect 68 700 102 733
rect 68 628 102 662
rect 68 556 102 590
rect 68 484 102 518
rect 68 412 102 446
rect 68 341 102 374
rect 68 340 100 341
rect 100 340 102 341
rect 68 270 102 302
rect 68 268 100 270
rect 100 268 102 270
rect 276 742 310 776
rect 348 742 356 776
rect 356 742 382 776
rect 420 742 424 776
rect 424 742 454 776
rect 492 742 526 776
rect 564 742 594 776
rect 594 742 598 776
rect 636 742 662 776
rect 662 742 670 776
rect 708 742 730 776
rect 730 742 742 776
rect 780 742 798 776
rect 798 742 814 776
rect 852 742 866 776
rect 866 742 886 776
rect 924 742 934 776
rect 934 742 958 776
rect 996 742 1030 776
rect 1068 742 1086 776
rect 1086 742 1102 776
rect 254 674 288 686
rect 254 652 288 674
rect 1086 662 1120 681
rect 475 626 490 660
rect 490 626 509 660
rect 547 626 558 660
rect 558 626 581 660
rect 619 626 626 660
rect 626 626 653 660
rect 691 626 694 660
rect 694 626 725 660
rect 763 626 796 660
rect 796 626 797 660
rect 835 626 864 660
rect 864 626 869 660
rect 907 626 932 660
rect 932 626 941 660
rect 979 626 1000 660
rect 1000 626 1013 660
rect 1086 647 1120 662
rect 254 572 288 604
rect 254 570 288 572
rect 254 504 288 522
rect 254 488 288 504
rect 254 436 288 441
rect 254 407 288 436
rect 336 565 370 572
rect 336 538 370 565
rect 336 497 370 500
rect 336 466 370 497
rect 1086 594 1120 609
rect 1086 575 1120 594
rect 1086 526 1120 537
rect 1086 503 1120 526
rect 1086 458 1120 465
rect 1086 431 1120 458
rect 474 370 490 404
rect 490 370 508 404
rect 556 370 558 404
rect 558 370 590 404
rect 637 370 660 404
rect 660 370 671 404
rect 718 370 728 404
rect 728 370 752 404
rect 799 370 830 404
rect 830 370 833 404
rect 880 370 898 404
rect 898 370 914 404
rect 961 370 966 404
rect 966 370 995 404
rect 1086 390 1120 393
rect 254 326 288 360
rect 1086 359 1120 390
rect 300 254 322 288
rect 322 254 334 288
rect 379 254 390 288
rect 390 254 413 288
rect 458 254 492 288
rect 537 254 560 288
rect 560 254 571 288
rect 616 254 628 288
rect 628 254 650 288
rect 695 254 696 288
rect 696 254 729 288
rect 774 254 798 288
rect 798 254 808 288
rect 852 254 866 288
rect 866 254 886 288
rect 930 254 934 288
rect 934 254 964 288
rect 1008 254 1042 288
rect 1086 254 1120 288
rect 1272 769 1306 803
rect 1272 697 1306 731
rect 1272 625 1306 659
rect 1272 554 1306 587
rect 1272 553 1306 554
rect 1272 483 1306 515
rect 1272 481 1306 483
rect 1272 412 1306 443
rect 1272 409 1306 412
rect 1272 341 1306 371
rect 1272 337 1306 341
rect 1272 270 1306 299
rect 1272 265 1306 270
rect 68 199 102 230
rect 68 196 100 199
rect 100 196 102 199
rect 68 124 102 158
rect 1272 198 1306 227
rect 1272 193 1306 198
rect 1272 126 1306 155
rect 1272 121 1306 126
rect 138 68 159 102
rect 159 68 172 102
rect 212 68 228 102
rect 228 68 246 102
rect 286 68 296 102
rect 296 68 320 102
rect 360 68 364 102
rect 364 68 394 102
rect 434 68 466 102
rect 466 68 468 102
rect 508 68 534 102
rect 534 68 542 102
rect 582 68 602 102
rect 602 68 616 102
rect 656 68 670 102
rect 670 68 690 102
rect 730 68 738 102
rect 738 68 764 102
rect 804 68 806 102
rect 806 68 838 102
rect 878 68 908 102
rect 908 68 912 102
rect 952 68 976 102
rect 976 68 986 102
rect 1026 68 1044 102
rect 1044 68 1060 102
rect 1100 68 1112 102
rect 1112 68 1134 102
rect 1174 68 1180 102
rect 1180 68 1208 102
<< metal1 >>
rect 1060 5355 1525 5380
rect 73 5239 79 5355
rect 195 5239 201 5355
rect 835 5239 841 5355
rect 1021 5239 1027 5355
rect 1060 5239 1066 5355
rect 1310 5239 1525 5355
rect 1060 5237 1525 5239
rect 1381 5178 1525 5237
rect 1507 5077 1525 5178
rect 385 4795 391 4911
rect 507 4795 513 4911
rect 1100 4795 1106 4911
rect 1222 4795 1228 4911
rect 1553 4795 1559 4911
rect 1675 4795 1681 4911
rect 582 4761 762 4767
rect 582 4639 762 4645
rect 1553 4611 1681 4795
rect 380 4495 386 4611
rect 502 4495 508 4611
rect 1100 4495 1106 4611
rect 1222 4495 1228 4611
rect 1553 4495 1559 4611
rect 1675 4495 1681 4611
rect 358 4339 536 4345
rect 358 3839 389 4339
rect 505 3839 536 4339
rect 358 3826 536 3839
rect 358 3774 389 3826
rect 441 3774 453 3826
rect 505 3774 536 3826
rect 358 3761 536 3774
rect 358 3709 389 3761
rect 441 3709 453 3761
rect 505 3709 536 3761
rect 358 3696 536 3709
rect 358 3644 389 3696
rect 441 3644 453 3696
rect 505 3644 536 3696
rect 358 3631 536 3644
rect 358 3579 389 3631
rect 441 3579 453 3631
rect 505 3579 536 3631
rect 1553 4229 1681 4495
rect 1553 3921 1559 4229
rect 1675 3998 1681 4229
rect 1675 3921 2051 3998
rect 1553 3908 2051 3921
rect 1553 3856 1559 3908
rect 1611 3856 1623 3908
rect 1675 3856 2051 3908
rect 1553 3778 2051 3856
rect 358 3566 536 3579
rect 358 3514 389 3566
rect 441 3514 453 3566
rect 505 3514 536 3566
rect 358 3501 536 3514
rect 358 3449 389 3501
rect 441 3449 453 3501
rect 505 3449 536 3501
rect 358 3443 536 3449
rect 66 3050 148 3249
rect 537 2927 669 2933
rect 537 2875 545 2927
rect 597 2875 609 2927
rect 661 2875 669 2927
rect 358 2861 536 2867
rect 358 2809 389 2861
rect 441 2809 453 2861
rect 505 2809 536 2861
rect 358 2796 536 2809
rect 358 2744 389 2796
rect 441 2744 453 2796
rect 505 2744 536 2796
rect 537 2828 669 2875
rect 537 2776 545 2828
rect 597 2776 609 2828
rect 661 2776 669 2828
rect 537 2770 669 2776
rect 358 2731 536 2744
rect 358 2679 389 2731
rect 441 2679 453 2731
rect 505 2679 536 2731
rect 358 2673 536 2679
rect 713 2673 719 3621
rect 835 2673 841 3621
rect 1444 3133 1470 3182
rect 886 2908 1088 2932
rect 886 2856 892 2908
rect 944 2856 961 2908
rect 1013 2856 1030 2908
rect 1082 2856 1088 2908
rect 886 2844 1088 2856
rect 886 2792 892 2844
rect 944 2792 961 2844
rect 1013 2792 1030 2844
rect 1082 2792 1088 2844
rect 886 2768 1088 2792
rect 1093 2861 1233 2867
rect 1093 2809 1105 2861
rect 1157 2809 1169 2861
rect 1221 2809 1233 2861
rect 1093 2796 1233 2809
rect 1093 2744 1105 2796
rect 1157 2744 1169 2796
rect 1221 2744 1233 2796
rect 1093 2731 1233 2744
rect 1093 2679 1105 2731
rect 1157 2679 1169 2731
rect 1221 2679 1233 2731
rect 1093 2673 1233 2679
rect 831 2611 1031 2617
rect 883 2559 905 2611
rect 957 2559 979 2611
rect 831 2517 1031 2559
rect 883 2465 905 2517
rect 957 2465 979 2517
rect 831 2459 1031 2465
rect 1553 2082 1681 3778
rect 1711 3121 1776 3237
rect 1892 3121 2113 3237
rect 385 1966 391 2082
rect 507 1966 513 2082
rect 572 2030 578 2082
rect 630 2030 646 2082
rect 698 2030 714 2082
rect 766 2030 772 2082
rect 572 2018 772 2030
rect 572 1966 578 2018
rect 630 1966 646 2018
rect 698 1966 714 2018
rect 766 1966 772 2018
rect 1104 1966 1110 2082
rect 1226 1966 1232 2082
rect 1553 1966 1559 2082
rect 1675 1966 1681 2082
rect 358 1189 514 1195
rect 410 1137 462 1189
rect 358 1090 514 1137
rect 410 1038 462 1090
rect 358 991 514 1038
rect 410 939 462 991
rect 358 933 514 939
rect 572 1189 772 1195
rect 624 1137 646 1189
rect 698 1137 720 1189
rect 572 1090 772 1137
rect 624 1038 646 1090
rect 698 1038 720 1090
rect 572 991 772 1038
rect 624 939 646 991
rect 698 939 720 991
rect 572 933 772 939
rect 831 1185 1031 1191
rect 883 1133 905 1185
rect 957 1133 979 1185
rect 831 1088 1031 1133
rect 883 1036 905 1088
rect 957 1036 979 1088
rect 831 991 1031 1036
rect 883 939 905 991
rect 957 939 979 991
rect 831 933 1031 939
tri 62 890 66 894 se
rect 66 890 108 933
tri 108 908 133 933 nw
tri 1228 908 1253 933 ne
rect 1253 908 1312 933
tri 1253 895 1266 908 ne
rect 62 878 108 890
rect 62 844 68 878
rect 102 844 108 878
rect 62 806 108 844
rect 62 772 68 806
rect 102 772 108 806
rect 62 734 108 772
rect 62 700 68 734
rect 102 700 108 734
rect 62 662 108 700
rect 62 628 68 662
rect 102 628 108 662
rect 62 590 108 628
rect 62 556 68 590
rect 102 556 108 590
rect 62 518 108 556
rect 62 484 68 518
rect 102 484 108 518
rect 62 446 108 484
rect 62 412 68 446
rect 102 412 108 446
rect 62 374 108 412
rect 62 340 68 374
rect 102 340 108 374
rect 62 302 108 340
rect 62 268 68 302
rect 102 268 108 302
rect 62 230 108 268
rect 248 825 364 877
rect 416 825 456 877
rect 508 825 578 877
rect 630 825 646 877
rect 698 825 714 877
rect 766 825 1132 877
rect 248 789 1132 825
rect 248 776 364 789
rect 416 776 456 789
rect 508 776 578 789
rect 630 776 646 789
rect 698 776 714 789
rect 766 776 1132 789
rect 248 742 276 776
rect 310 742 348 776
rect 416 742 420 776
rect 454 742 456 776
rect 526 742 564 776
rect 630 742 636 776
rect 698 742 708 776
rect 766 742 780 776
rect 814 742 852 776
rect 886 742 924 776
rect 958 742 996 776
rect 1030 742 1068 776
rect 1102 742 1132 776
rect 248 737 364 742
rect 416 737 456 742
rect 508 737 578 742
rect 630 737 646 742
rect 698 737 714 742
rect 766 737 1132 742
rect 248 736 1132 737
rect 248 731 327 736
tri 327 731 332 736 nw
tri 1042 731 1047 736 ne
rect 1047 731 1132 736
rect 248 686 294 731
tri 294 698 327 731 nw
tri 1047 698 1080 731 ne
rect 248 652 254 686
rect 288 652 294 686
rect 1080 681 1132 731
rect 248 604 294 652
rect 463 660 650 669
rect 702 660 714 669
rect 766 660 778 669
rect 830 660 842 669
rect 463 626 475 660
rect 509 626 547 660
rect 581 626 619 660
rect 830 626 835 660
rect 463 617 650 626
rect 702 617 714 626
rect 766 617 778 626
rect 830 617 842 626
rect 894 617 906 669
rect 958 617 970 669
rect 1022 617 1028 669
rect 1080 647 1086 681
rect 1120 647 1132 681
rect 248 570 254 604
rect 288 570 294 604
rect 1080 609 1132 647
rect 248 522 294 570
rect 248 488 254 522
rect 288 488 294 522
rect 248 441 294 488
rect 327 577 379 584
rect 327 513 379 525
rect 327 454 379 461
rect 1080 575 1086 609
rect 1120 575 1132 609
rect 1080 537 1132 575
rect 1080 503 1086 537
rect 1120 503 1132 537
rect 1080 465 1132 503
rect 248 407 254 441
rect 288 407 294 441
rect 1080 431 1086 465
rect 1120 431 1132 465
rect 248 360 294 407
rect 462 404 837 413
rect 889 404 901 413
rect 953 404 1007 413
rect 462 370 474 404
rect 508 370 556 404
rect 590 370 637 404
rect 671 370 718 404
rect 752 370 799 404
rect 833 370 837 404
rect 953 370 961 404
rect 995 370 1007 404
rect 462 361 837 370
rect 889 361 901 370
rect 953 361 1007 370
rect 1080 393 1132 431
rect 248 326 254 360
rect 288 326 294 360
rect 1080 359 1086 393
rect 1120 359 1132 393
rect 248 314 294 326
tri 294 314 312 332 sw
tri 1062 314 1080 332 se
rect 1080 314 1132 359
rect 248 299 312 314
tri 312 299 327 314 sw
tri 1047 299 1062 314 se
rect 1062 299 1132 314
rect 248 294 327 299
tri 327 294 332 299 sw
tri 1042 294 1047 299 se
rect 1047 294 1132 299
rect 248 288 1132 294
rect 248 254 300 288
rect 334 254 379 288
rect 413 254 458 288
rect 492 254 537 288
rect 571 254 616 288
rect 650 254 695 288
rect 729 254 774 288
rect 808 254 852 288
rect 886 254 930 288
rect 964 254 1008 288
rect 1042 254 1086 288
rect 1120 254 1132 288
rect 248 242 1132 254
rect 1266 875 1312 908
tri 1312 895 1350 933 nw
rect 1266 841 1272 875
rect 1306 841 1312 875
rect 1865 851 1967 853
rect 1266 803 1312 841
rect 1711 828 2113 851
rect 1266 769 1272 803
rect 1306 769 1312 803
rect 1266 731 1312 769
rect 1266 697 1272 731
rect 1306 697 1312 731
rect 1266 659 1312 697
rect 1266 625 1272 659
rect 1306 625 1312 659
rect 1266 587 1312 625
rect 1266 553 1272 587
rect 1306 553 1312 587
rect 1266 515 1312 553
rect 1266 481 1272 515
rect 1306 481 1312 515
rect 1266 443 1312 481
rect 1266 409 1272 443
rect 1306 409 1312 443
rect 1266 371 1312 409
rect 1266 337 1272 371
rect 1306 337 1312 371
rect 1266 299 1312 337
rect 1266 265 1272 299
rect 1306 265 1312 299
rect 62 196 68 230
rect 102 196 108 230
rect 62 158 108 196
rect 62 124 68 158
rect 102 124 108 158
rect 1266 227 1312 265
rect 1266 193 1272 227
rect 1306 193 1312 227
rect 1266 155 1312 193
rect 62 121 108 124
tri 108 121 133 146 sw
tri 1255 135 1266 146 se
rect 1266 135 1272 155
tri 1241 121 1255 135 se
rect 1255 121 1272 135
rect 1306 121 1312 155
rect 62 108 133 121
tri 133 108 146 121 sw
tri 1228 108 1241 121 se
rect 1241 108 1312 121
rect 62 102 1312 108
rect 62 68 138 102
rect 172 68 212 102
rect 246 68 286 102
rect 320 68 360 102
rect 394 68 434 102
rect 468 68 508 102
rect 542 68 582 102
rect 616 68 656 102
rect 690 68 730 102
rect 764 68 804 102
rect 838 68 878 102
rect 912 68 952 102
rect 986 68 1026 102
rect 1060 68 1100 102
rect 1134 68 1174 102
rect 1208 68 1312 102
rect 62 56 1312 68
<< via1 >>
rect 79 5239 195 5355
rect 841 5335 1021 5355
rect 841 5301 843 5335
rect 843 5301 877 5335
rect 877 5301 915 5335
rect 915 5301 949 5335
rect 949 5301 987 5335
rect 987 5301 1021 5335
rect 841 5239 1021 5301
rect 1066 5239 1310 5355
rect 391 4795 507 4911
rect 1106 4795 1222 4911
rect 1559 4795 1675 4911
rect 582 4645 762 4761
rect 386 4495 502 4611
rect 1106 4495 1222 4611
rect 1559 4495 1675 4611
rect 389 3839 505 4339
rect 389 3774 441 3826
rect 453 3774 505 3826
rect 389 3709 441 3761
rect 453 3709 505 3761
rect 389 3644 441 3696
rect 453 3644 505 3696
rect 389 3579 441 3631
rect 453 3579 505 3631
rect 1559 3921 1675 4229
rect 1559 3856 1611 3908
rect 1623 3856 1675 3908
rect 389 3514 441 3566
rect 453 3514 505 3566
rect 389 3449 441 3501
rect 453 3449 505 3501
rect 545 2875 597 2927
rect 609 2875 661 2927
rect 389 2809 441 2861
rect 453 2809 505 2861
rect 389 2744 441 2796
rect 453 2744 505 2796
rect 545 2776 597 2828
rect 609 2776 661 2828
rect 389 2679 441 2731
rect 453 2679 505 2731
rect 719 2673 835 3621
rect 892 2856 944 2908
rect 961 2856 1013 2908
rect 1030 2856 1082 2908
rect 892 2792 944 2844
rect 961 2792 1013 2844
rect 1030 2792 1082 2844
rect 1105 2809 1157 2861
rect 1169 2809 1221 2861
rect 1105 2744 1157 2796
rect 1169 2744 1221 2796
rect 1105 2679 1157 2731
rect 1169 2679 1221 2731
rect 831 2559 883 2611
rect 905 2559 957 2611
rect 979 2559 1031 2611
rect 831 2465 883 2517
rect 905 2465 957 2517
rect 979 2465 1031 2517
rect 1776 3121 1892 3237
rect 391 1966 507 2082
rect 578 2030 630 2082
rect 646 2030 698 2082
rect 714 2030 766 2082
rect 578 1966 630 2018
rect 646 1966 698 2018
rect 714 1966 766 2018
rect 1110 1966 1226 2082
rect 1559 1966 1675 2082
rect 358 1137 410 1189
rect 462 1137 514 1189
rect 358 1038 410 1090
rect 462 1038 514 1090
rect 358 939 410 991
rect 462 939 514 991
rect 572 1137 624 1189
rect 646 1137 698 1189
rect 720 1137 772 1189
rect 572 1038 624 1090
rect 646 1038 698 1090
rect 720 1038 772 1090
rect 572 939 624 991
rect 646 939 698 991
rect 720 939 772 991
rect 831 1133 883 1185
rect 905 1133 957 1185
rect 979 1133 1031 1185
rect 831 1036 883 1088
rect 905 1036 957 1088
rect 979 1036 1031 1088
rect 831 939 883 991
rect 905 939 957 991
rect 979 939 1031 991
rect 364 825 416 877
rect 456 825 508 877
rect 578 825 630 877
rect 646 825 698 877
rect 714 825 766 877
rect 364 776 416 789
rect 456 776 508 789
rect 578 776 630 789
rect 646 776 698 789
rect 714 776 766 789
rect 364 742 382 776
rect 382 742 416 776
rect 456 742 492 776
rect 492 742 508 776
rect 578 742 598 776
rect 598 742 630 776
rect 646 742 670 776
rect 670 742 698 776
rect 714 742 742 776
rect 742 742 766 776
rect 364 737 416 742
rect 456 737 508 742
rect 578 737 630 742
rect 646 737 698 742
rect 714 737 766 742
rect 650 660 702 669
rect 714 660 766 669
rect 778 660 830 669
rect 842 660 894 669
rect 650 626 653 660
rect 653 626 691 660
rect 691 626 702 660
rect 714 626 725 660
rect 725 626 763 660
rect 763 626 766 660
rect 778 626 797 660
rect 797 626 830 660
rect 842 626 869 660
rect 869 626 894 660
rect 650 617 702 626
rect 714 617 766 626
rect 778 617 830 626
rect 842 617 894 626
rect 906 660 958 669
rect 906 626 907 660
rect 907 626 941 660
rect 941 626 958 660
rect 906 617 958 626
rect 970 660 1022 669
rect 970 626 979 660
rect 979 626 1013 660
rect 1013 626 1022 660
rect 970 617 1022 626
rect 327 572 379 577
rect 327 538 336 572
rect 336 538 370 572
rect 370 538 379 572
rect 327 525 379 538
rect 327 500 379 513
rect 327 466 336 500
rect 336 466 370 500
rect 370 466 379 500
rect 327 461 379 466
rect 837 404 889 413
rect 901 404 953 413
rect 837 370 880 404
rect 880 370 889 404
rect 901 370 914 404
rect 914 370 953 404
rect 837 361 889 370
rect 901 361 953 370
<< metal2 >>
rect 0 5239 79 5355
rect 195 5239 841 5355
rect 1021 5239 1066 5355
rect 1310 5239 1316 5355
rect 358 4795 391 4911
rect 507 4795 1106 4911
rect 1222 4795 1559 4911
rect 1675 4795 1681 4911
rect 358 4761 1898 4767
rect 358 4645 582 4761
rect 762 4645 1898 4761
rect 358 4639 1898 4645
tri 1736 4611 1764 4639 ne
rect 1764 4611 1898 4639
rect 358 4495 386 4611
rect 502 4495 1106 4611
rect 1222 4495 1559 4611
rect 1675 4495 1681 4611
tri 1764 4605 1770 4611 ne
rect 358 4339 1233 4345
rect 358 3839 389 4339
rect 505 3839 1233 4339
rect 358 3826 1233 3839
rect 358 3774 389 3826
rect 441 3774 453 3826
rect 505 3774 1233 3826
rect 358 3761 1233 3774
rect 358 3709 389 3761
rect 441 3709 453 3761
rect 505 3709 1233 3761
rect 358 3696 1233 3709
rect 358 3644 389 3696
rect 441 3644 453 3696
rect 505 3644 1233 3696
rect 358 3631 1233 3644
rect 358 3579 389 3631
rect 441 3579 453 3631
rect 505 3621 1233 3631
rect 505 3579 719 3621
rect 358 3566 719 3579
rect 358 3514 389 3566
rect 441 3514 453 3566
rect 505 3514 719 3566
rect 358 3501 719 3514
rect 358 3449 389 3501
rect 441 3449 453 3501
rect 505 3449 719 3501
rect 358 2927 719 3449
rect 358 2875 545 2927
rect 597 2875 609 2927
rect 661 2875 719 2927
rect 358 2861 719 2875
rect 358 2809 389 2861
rect 441 2809 453 2861
rect 505 2828 719 2861
rect 505 2809 545 2828
rect 358 2796 545 2809
rect 358 2744 389 2796
rect 441 2744 453 2796
rect 505 2776 545 2796
rect 597 2776 609 2828
rect 661 2776 719 2828
rect 505 2744 719 2776
rect 358 2731 719 2744
rect 358 2679 389 2731
rect 441 2679 453 2731
rect 505 2679 719 2731
rect 358 2673 719 2679
rect 835 3121 1233 3621
rect 1553 4229 1681 4235
rect 1553 3921 1559 4229
rect 1675 3921 1681 4229
rect 1553 3908 1681 3921
rect 1553 3856 1559 3908
rect 1611 3856 1623 3908
rect 1675 3856 1681 3908
tri 1233 3121 1299 3187 sw
rect 835 3015 1299 3121
tri 1299 3015 1405 3121 sw
rect 835 2981 1405 3015
tri 1405 2981 1439 3015 sw
tri 1519 2981 1553 3015 se
rect 1553 2981 1681 3856
rect 835 2908 1681 2981
rect 835 2856 892 2908
rect 944 2856 961 2908
rect 1013 2856 1030 2908
rect 1082 2861 1681 2908
rect 1082 2856 1105 2861
rect 835 2844 1105 2856
rect 835 2792 892 2844
rect 944 2792 961 2844
rect 1013 2792 1030 2844
rect 1082 2809 1105 2844
rect 1157 2809 1169 2861
rect 1221 2809 1681 2861
rect 1082 2796 1681 2809
rect 1082 2792 1105 2796
rect 835 2744 1105 2792
rect 1157 2744 1169 2796
rect 1221 2744 1681 2796
rect 835 2731 1681 2744
rect 835 2679 1105 2731
rect 1157 2679 1169 2731
rect 1221 2679 1681 2731
rect 835 2673 1681 2679
rect 1770 3237 1898 4611
rect 1770 3121 1776 3237
rect 1892 3121 1898 3237
tri 1736 2617 1770 2651 se
rect 1770 2617 1898 3121
rect 822 2611 1898 2617
rect 822 2559 831 2611
rect 883 2559 905 2611
rect 957 2559 979 2611
rect 1031 2559 1898 2611
rect 822 2517 1898 2559
rect 822 2465 831 2517
rect 883 2465 905 2517
rect 957 2465 979 2517
rect 1031 2465 1898 2517
rect 822 2459 1898 2465
rect 358 1966 391 2082
rect 507 2030 578 2082
rect 630 2030 646 2082
rect 698 2030 714 2082
rect 766 2030 1110 2082
rect 507 2018 1110 2030
rect 507 1966 578 2018
rect 630 1966 646 2018
rect 698 1966 714 2018
rect 766 1966 1110 2018
rect 1226 1966 1559 2082
rect 1675 1966 1681 2082
rect 358 1189 514 1195
rect 410 1137 462 1189
rect 358 1090 514 1137
rect 410 1038 462 1090
rect 358 991 514 1038
rect 410 939 462 991
rect 358 877 514 939
rect 358 825 364 877
rect 416 825 456 877
rect 508 825 514 877
rect 358 789 514 825
rect 358 737 364 789
rect 416 737 456 789
rect 508 737 514 789
rect 358 736 514 737
rect 572 1189 772 1195
rect 624 1137 646 1189
rect 698 1137 720 1189
rect 572 1090 772 1137
rect 624 1038 646 1090
rect 698 1038 720 1090
rect 572 991 772 1038
rect 624 939 646 991
rect 698 939 720 991
rect 572 877 772 939
rect 572 825 578 877
rect 630 825 646 877
rect 698 825 714 877
rect 766 825 772 877
rect 572 789 772 825
rect 572 737 578 789
rect 630 737 646 789
rect 698 737 714 789
rect 766 737 772 789
rect 572 736 772 737
rect 831 1185 1031 1191
rect 883 1133 905 1185
rect 957 1133 979 1185
rect 831 1088 1031 1133
rect 883 1036 905 1088
rect 957 1036 979 1088
rect 831 991 1031 1036
rect 883 939 905 991
rect 957 939 979 991
tri 793 669 831 707 se
rect 831 669 1031 939
rect 644 617 650 669
rect 702 617 714 669
rect 766 617 778 669
rect 830 617 842 669
rect 894 617 906 669
rect 958 617 970 669
rect 1022 617 1031 669
rect 327 577 1483 583
rect 379 525 1483 577
rect 327 513 1483 525
rect 379 461 1483 513
rect 327 455 1483 461
rect 831 361 837 413
rect 889 361 901 413
rect 953 361 1478 413
use sky130_fd_io__res250only_small  sky130_fd_io__res250only_small_0
timestamp 1683767628
transform 0 -1 2114 1 0 851
box 0 0 2270 404
use sky130_fd_io__signal_5_sym_hv_local_5term  sky130_fd_io__signal_5_sym_hv_local_5term_0
timestamp 1683767628
transform 1 0 0 0 1 867
box 0 0 1591 2424
use sky130_fd_io__signal_5_sym_hv_local_5term  sky130_fd_io__signal_5_sym_hv_local_5term_1
timestamp 1683767628
transform 1 0 0 0 -1 5443
box 0 0 1591 2424
use sky130_fd_pr__nfet_01v8__example_55959141808555  sky130_fd_pr__nfet_01v8__example_55959141808555_0
timestamp 1683767628
transform 0 -1 1012 1 0 415
box -1 0 201 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1683767628
transform 0 -1 370 -1 0 572
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_0
timestamp 1683767628
transform 0 1 843 -1 0 5335
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808290  sky130_fd_pr__via_l1m1__example_55959141808290_0
timestamp 1683767628
transform 1 0 475 0 -1 660
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808326  sky130_fd_pr__via_l1m1__example_55959141808326_0
timestamp 1683767628
transform 0 -1 102 1 0 124
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808326  sky130_fd_pr__via_l1m1__example_55959141808326_1
timestamp 1683767628
transform 0 -1 1306 -1 0 875
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808372  sky130_fd_pr__via_l1m1__example_55959141808372_0
timestamp 1683767628
transform 0 -1 1120 -1 0 681
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808400  sky130_fd_pr__via_l1m1__example_55959141808400_0
timestamp 1683767628
transform 1 0 276 0 1 742
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1683767628
transform 0 -1 379 1 0 455
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_0
timestamp 1683767628
transform 1 0 73 0 1 5239
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_1
timestamp 1683767628
transform -1 0 1232 0 -1 2082
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_2
timestamp 1683767628
transform 1 0 385 0 -1 4911
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_3
timestamp 1683767628
transform 1 0 1100 0 -1 4611
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_4
timestamp 1683767628
transform 1 0 1100 0 1 4795
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_5
timestamp 1683767628
transform 1 0 385 0 -1 2082
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_6
timestamp 1683767628
transform 1 0 1553 0 -1 2082
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_7
timestamp 1683767628
transform 1 0 380 0 -1 4611
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808402  sky130_fd_pr__via_m1m2__example_55959141808402_0
timestamp 1683767628
transform 0 1 582 1 0 4639
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808551  sky130_fd_pr__via_m1m2__example_55959141808551_0
timestamp 1683767628
transform -1 0 1316 0 1 5239
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808552  sky130_fd_pr__via_m1m2__example_55959141808552_0
timestamp 1683767628
transform 1 0 835 0 1 5239
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808553  sky130_fd_pr__via_m1m2__example_55959141808553_0
timestamp 1683767628
transform -1 0 1028 0 -1 669
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808554  sky130_fd_pr__via_m1m2__example_55959141808554_0
timestamp 1683767628
transform 1 0 713 0 1 2673
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_0
timestamp 1683767628
transform -1 0 386 0 -1 615
box 0 0 1 1
<< labels >>
flabel metal2 s 1375 370 1474 407 3 FreeSans 200 0 0 0 OUT_VT
port 2 nsew
flabel metal2 s 1375 469 1469 567 3 FreeSans 200 0 0 0 VTRIP_SEL_H
port 3 nsew
flabel metal2 s 88 5277 260 5345 3 FreeSans 520 0 0 0 VDDIO_Q
port 1 nsew
flabel metal1 s 1865 831 1967 853 3 FreeSans 520 0 0 0 IN_H
port 5 nsew
flabel metal1 s 2074 3125 2113 3234 7 FreeSans 200 0 0 0 OUT_H
port 6 nsew
flabel metal1 s 1700 3778 2042 3994 3 FreeSans 200 0 0 0 VSSD
port 7 nsew
<< properties >>
string GDS_END 35964742
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 35939170
<< end >>
