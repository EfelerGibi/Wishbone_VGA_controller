magic
tech sky130A
timestamp 1683767628
<< properties >>
string GDS_END 37308604
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 37306488
<< end >>
