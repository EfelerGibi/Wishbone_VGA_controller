magic
tech sky130B
magscale 1 2
timestamp 1683767628
<< pwell >>
rect 467 350 491 401
<< obsli1 >>
rect 0 852 876 918
rect 0 746 66 852
rect 100 782 776 816
rect 0 712 377 746
rect 0 606 66 712
rect 411 676 465 782
rect 810 746 876 852
rect 499 712 876 746
rect 100 642 776 676
rect 0 572 377 606
rect 0 346 66 572
rect 411 536 465 642
rect 810 606 876 712
rect 499 572 876 606
rect 100 502 776 536
rect 411 416 465 502
rect 100 382 776 416
rect 0 312 377 346
rect 0 206 66 312
rect 411 276 465 382
rect 810 346 876 572
rect 499 312 876 346
rect 100 242 776 276
rect 0 172 377 206
rect 0 66 66 172
rect 411 136 465 242
rect 810 206 876 312
rect 499 172 876 206
rect 100 102 776 136
rect 810 66 876 172
rect 0 0 876 66
<< obsm1 >>
rect 0 852 876 918
rect 0 66 66 852
rect 113 491 141 824
rect 169 519 197 852
rect 225 491 253 824
rect 281 519 309 852
rect 337 491 365 824
rect 411 491 465 824
rect 511 491 539 824
rect 567 519 595 852
rect 623 491 651 824
rect 679 519 707 852
rect 735 491 763 824
rect 113 427 763 491
rect 113 94 141 427
rect 169 66 197 399
rect 225 94 253 427
rect 281 66 309 399
rect 337 94 365 427
rect 411 94 465 427
rect 511 94 539 427
rect 567 66 595 399
rect 623 94 651 427
rect 679 66 707 399
rect 735 94 763 427
rect 810 66 876 852
rect 0 0 876 66
<< metal2 >>
rect 0 852 383 918
rect 0 768 66 852
rect 411 824 465 918
rect 493 852 876 918
rect 94 796 782 824
rect 0 740 383 768
rect 0 656 66 740
rect 411 712 465 796
rect 810 768 876 852
rect 493 740 876 768
rect 94 684 782 712
rect 0 628 383 656
rect 0 544 66 628
rect 411 600 465 684
rect 810 656 876 740
rect 493 628 876 656
rect 94 572 782 600
rect 0 516 383 544
rect 0 514 66 516
rect 411 486 465 572
rect 810 544 876 628
rect 493 516 876 544
rect 810 514 876 516
rect 0 432 876 486
rect 0 402 66 404
rect 0 374 383 402
rect 0 290 66 374
rect 411 346 465 432
rect 810 402 876 404
rect 493 374 876 402
rect 94 318 782 346
rect 0 262 383 290
rect 0 178 66 262
rect 411 234 465 318
rect 810 290 876 374
rect 493 262 876 290
rect 94 206 782 234
rect 0 150 383 178
rect 0 66 66 150
rect 411 122 465 206
rect 810 178 876 262
rect 493 150 876 178
rect 94 94 782 122
rect 0 0 383 66
rect 411 0 465 94
rect 810 66 876 150
rect 493 0 876 66
<< metal3 >>
rect 0 0 876 918
<< labels >>
rlabel metal2 s 810 768 876 852 6 C0
port 1 nsew
rlabel metal2 s 810 656 876 740 6 C0
port 1 nsew
rlabel metal2 s 810 544 876 628 6 C0
port 1 nsew
rlabel metal2 s 810 514 876 516 6 C0
port 1 nsew
rlabel metal2 s 810 402 876 404 6 C0
port 1 nsew
rlabel metal2 s 810 290 876 374 6 C0
port 1 nsew
rlabel metal2 s 810 178 876 262 6 C0
port 1 nsew
rlabel metal2 s 810 66 876 150 6 C0
port 1 nsew
rlabel metal2 s 493 852 876 918 6 C0
port 1 nsew
rlabel metal2 s 493 740 876 768 6 C0
port 1 nsew
rlabel metal2 s 493 628 876 656 6 C0
port 1 nsew
rlabel metal2 s 493 516 876 544 6 C0
port 1 nsew
rlabel metal2 s 493 374 876 402 6 C0
port 1 nsew
rlabel metal2 s 493 262 876 290 6 C0
port 1 nsew
rlabel metal2 s 493 150 876 178 6 C0
port 1 nsew
rlabel metal2 s 493 0 876 66 6 C0
port 1 nsew
rlabel metal2 s 0 852 383 918 6 C0
port 1 nsew
rlabel metal2 s 0 768 66 852 6 C0
port 1 nsew
rlabel metal2 s 0 740 383 768 6 C0
port 1 nsew
rlabel metal2 s 0 656 66 740 6 C0
port 1 nsew
rlabel metal2 s 0 628 383 656 6 C0
port 1 nsew
rlabel metal2 s 0 544 66 628 6 C0
port 1 nsew
rlabel metal2 s 0 516 383 544 6 C0
port 1 nsew
rlabel metal2 s 0 514 66 516 6 C0
port 1 nsew
rlabel metal2 s 0 402 66 404 6 C0
port 1 nsew
rlabel metal2 s 0 374 383 402 6 C0
port 1 nsew
rlabel metal2 s 0 290 66 374 6 C0
port 1 nsew
rlabel metal2 s 0 262 383 290 6 C0
port 1 nsew
rlabel metal2 s 0 178 66 262 6 C0
port 1 nsew
rlabel metal2 s 0 150 383 178 6 C0
port 1 nsew
rlabel metal2 s 0 66 66 150 6 C0
port 1 nsew
rlabel metal2 s 0 0 383 66 6 C0
port 1 nsew
rlabel metal2 s 411 824 465 918 6 C1
port 2 nsew
rlabel metal2 s 411 712 465 796 6 C1
port 2 nsew
rlabel metal2 s 411 600 465 684 6 C1
port 2 nsew
rlabel metal2 s 411 486 465 572 6 C1
port 2 nsew
rlabel metal2 s 411 346 465 432 6 C1
port 2 nsew
rlabel metal2 s 411 234 465 318 6 C1
port 2 nsew
rlabel metal2 s 411 122 465 206 6 C1
port 2 nsew
rlabel metal2 s 411 0 465 94 6 C1
port 2 nsew
rlabel metal2 s 94 796 782 824 6 C1
port 2 nsew
rlabel metal2 s 94 684 782 712 6 C1
port 2 nsew
rlabel metal2 s 94 572 782 600 6 C1
port 2 nsew
rlabel metal2 s 94 318 782 346 6 C1
port 2 nsew
rlabel metal2 s 94 206 782 234 6 C1
port 2 nsew
rlabel metal2 s 94 94 782 122 6 C1
port 2 nsew
rlabel metal2 s 0 432 876 486 6 C1
port 2 nsew
rlabel metal3 s 0 0 876 918 6 MET3
port 4 nsew
rlabel pwell s 467 350 491 401 6 SUB
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 876 918
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 99422
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 81886
string device primitive
<< end >>
