magic
tech sky130A
magscale 1 2
timestamp 1683767628
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 1 145 541 157
rect 825 145 1103 203
rect 1 21 1103 145
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 435 47 465 131
rect 530 47 560 119
rect 629 47 659 119
rect 713 47 743 119
rect 903 47 933 177
rect 990 47 1020 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 369 381 497
rect 435 369 465 497
rect 530 413 560 497
rect 614 413 644 497
rect 713 413 743 497
rect 903 297 933 497
rect 990 297 1020 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 119 351 131
rect 299 85 307 119
rect 341 85 351 119
rect 299 47 351 85
rect 381 89 435 131
rect 381 55 391 89
rect 425 55 435 89
rect 381 47 435 55
rect 465 119 515 131
rect 851 133 903 177
rect 465 47 530 119
rect 560 107 629 119
rect 560 73 584 107
rect 618 73 629 107
rect 560 47 629 73
rect 659 47 713 119
rect 743 106 795 119
rect 743 72 753 106
rect 787 72 795 106
rect 743 47 795 72
rect 851 99 859 133
rect 893 99 903 133
rect 851 47 903 99
rect 933 127 990 177
rect 933 93 946 127
rect 980 93 990 127
rect 933 47 990 93
rect 1020 133 1077 177
rect 1020 99 1035 133
rect 1069 99 1077 133
rect 1020 47 1077 99
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 483 351 497
rect 299 449 307 483
rect 341 449 351 483
rect 299 415 351 449
rect 299 381 307 415
rect 341 381 351 415
rect 299 369 351 381
rect 381 485 435 497
rect 381 451 391 485
rect 425 451 435 485
rect 381 417 435 451
rect 381 383 391 417
rect 425 383 435 417
rect 381 369 435 383
rect 465 413 530 497
rect 560 485 614 497
rect 560 451 570 485
rect 604 451 614 485
rect 560 413 614 451
rect 644 413 713 497
rect 743 477 797 497
rect 743 443 755 477
rect 789 443 797 477
rect 743 413 797 443
rect 851 471 903 497
rect 851 437 859 471
rect 893 437 903 471
rect 465 369 515 413
rect 851 368 903 437
rect 851 334 859 368
rect 893 334 903 368
rect 851 297 903 334
rect 933 484 990 497
rect 933 450 946 484
rect 980 450 990 484
rect 933 364 990 450
rect 933 330 946 364
rect 980 330 990 364
rect 933 297 990 330
rect 1020 475 1077 497
rect 1020 441 1035 475
rect 1069 441 1077 475
rect 1020 384 1077 441
rect 1020 350 1035 384
rect 1069 350 1077 384
rect 1020 297 1077 350
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 85 341 119
rect 391 55 425 89
rect 584 73 618 107
rect 753 72 787 106
rect 859 99 893 133
rect 946 93 980 127
rect 1035 99 1069 133
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 449 341 483
rect 307 381 341 415
rect 391 451 425 485
rect 391 383 425 417
rect 570 451 604 485
rect 755 443 789 477
rect 859 437 893 471
rect 859 334 893 368
rect 946 450 980 484
rect 946 330 980 364
rect 1035 441 1069 475
rect 1035 350 1069 384
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 435 497 465 523
rect 530 497 560 523
rect 614 497 644 523
rect 713 497 743 523
rect 903 497 933 523
rect 990 497 1020 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 280 76 318
rect 22 264 76 280
rect 163 274 193 363
rect 22 230 32 264
rect 66 230 76 264
rect 22 214 76 230
rect 118 264 193 274
rect 118 230 134 264
rect 168 230 193 264
rect 351 241 381 369
rect 118 220 193 230
rect 46 176 76 214
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 298 225 381 241
rect 298 191 308 225
rect 342 191 381 225
rect 435 219 465 369
rect 530 337 560 413
rect 614 375 644 413
rect 603 365 669 375
rect 507 321 561 337
rect 603 331 619 365
rect 653 331 669 365
rect 603 321 669 331
rect 713 373 743 413
rect 713 357 812 373
rect 713 323 768 357
rect 802 323 812 357
rect 507 287 517 321
rect 551 287 561 321
rect 507 279 561 287
rect 713 307 812 323
rect 507 271 659 279
rect 531 249 659 271
rect 298 175 381 191
rect 351 131 381 175
rect 424 203 478 219
rect 424 169 434 203
rect 468 169 478 203
rect 424 153 478 169
rect 530 191 587 207
rect 530 157 543 191
rect 577 157 587 191
rect 435 131 465 153
rect 530 141 587 157
rect 530 119 560 141
rect 629 119 659 249
rect 713 119 743 307
rect 903 265 933 297
rect 990 265 1020 297
rect 791 249 933 265
rect 791 215 801 249
rect 835 215 933 249
rect 791 199 933 215
rect 975 249 1029 265
rect 975 215 985 249
rect 1019 215 1029 249
rect 975 199 1029 215
rect 903 177 933 199
rect 990 177 1020 199
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 435 21 465 47
rect 530 21 560 47
rect 629 21 659 47
rect 713 21 743 47
rect 903 21 933 47
rect 990 21 1020 47
<< polycont >>
rect 32 230 66 264
rect 134 230 168 264
rect 308 191 342 225
rect 619 331 653 365
rect 768 323 802 357
rect 517 287 551 321
rect 434 169 468 203
rect 543 157 577 191
rect 801 215 835 249
rect 985 215 1019 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 391 485 454 527
rect 237 443 248 477
rect 203 409 248 443
rect 69 375 156 393
rect 35 359 156 375
rect 18 264 66 325
rect 18 230 32 264
rect 18 197 66 230
rect 122 323 156 359
rect 122 280 156 289
rect 237 391 248 409
rect 203 357 214 375
rect 203 337 248 357
rect 291 449 307 483
rect 341 449 357 483
rect 291 415 357 449
rect 291 381 307 415
rect 341 381 357 415
rect 122 264 168 280
rect 122 230 134 264
rect 122 214 168 230
rect 122 161 156 214
rect 35 127 156 161
rect 35 119 69 127
rect 203 119 237 337
rect 291 333 357 381
rect 425 451 454 485
rect 554 451 570 485
rect 604 451 721 485
rect 391 417 454 451
rect 425 383 454 417
rect 391 367 454 383
rect 585 391 653 399
rect 585 357 586 391
rect 620 365 653 391
rect 291 299 428 333
rect 292 225 358 265
rect 292 191 308 225
rect 342 191 358 225
rect 394 219 428 299
rect 494 323 551 337
rect 528 321 551 323
rect 494 287 517 289
rect 494 271 551 287
rect 585 331 619 357
rect 585 315 653 331
rect 394 203 468 219
rect 585 207 619 315
rect 687 265 721 451
rect 755 477 789 527
rect 755 427 789 443
rect 859 471 903 487
rect 893 437 903 471
rect 859 373 903 437
rect 768 368 903 373
rect 768 357 859 368
rect 802 334 859 357
rect 893 334 903 368
rect 802 323 903 334
rect 768 307 903 323
rect 939 484 980 527
rect 939 450 946 484
rect 939 364 980 450
rect 939 330 946 364
rect 1030 475 1087 491
rect 1030 441 1035 475
rect 1069 441 1087 475
rect 1030 384 1087 441
rect 1030 350 1035 384
rect 1069 350 1087 384
rect 1030 334 1087 350
rect 939 314 980 330
rect 869 265 903 307
rect 687 249 835 265
rect 687 233 801 249
rect 394 169 434 203
rect 394 157 468 169
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 203 69 237 85
rect 307 153 468 157
rect 543 191 619 207
rect 577 157 619 191
rect 307 123 428 153
rect 543 141 619 157
rect 666 215 801 233
rect 666 199 835 215
rect 869 249 1019 265
rect 869 215 985 249
rect 869 199 1019 215
rect 307 119 341 123
rect 666 107 700 199
rect 869 149 903 199
rect 1053 149 1087 334
rect 307 69 341 85
rect 103 17 169 59
rect 375 55 391 89
rect 425 55 441 89
rect 568 73 584 107
rect 618 73 700 107
rect 859 133 903 149
rect 375 17 441 55
rect 737 72 753 106
rect 787 72 803 106
rect 893 99 903 133
rect 859 83 903 99
rect 939 127 980 143
rect 939 93 946 127
rect 737 17 803 72
rect 939 17 980 93
rect 1030 133 1087 149
rect 1030 99 1035 133
rect 1069 99 1087 133
rect 1030 83 1087 99
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 122 289 156 323
rect 214 375 237 391
rect 237 375 248 391
rect 214 357 248 375
rect 586 365 620 391
rect 586 357 619 365
rect 619 357 620 365
rect 494 321 528 323
rect 494 289 517 321
rect 517 289 528 321
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 574 391 632 397
rect 574 388 586 391
rect 248 360 586 388
rect 248 357 260 360
rect 202 351 260 357
rect 574 357 586 360
rect 620 357 632 391
rect 574 351 632 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 482 323 540 329
rect 482 320 494 323
rect 156 292 494 320
rect 156 289 168 292
rect 110 283 168 289
rect 482 289 494 292
rect 528 289 540 323
rect 482 283 540 289
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel locali s 310 221 344 255 0 FreeSans 200 0 0 0 D
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1046 357 1080 391 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1046 425 1080 459 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 1046 85 1080 119 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
rlabel comment s 0 0 0 0 4 dlxtp_1
rlabel metal1 s 0 -48 1104 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1104 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_END 2892046
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2881896
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 27.600 0.000 
<< end >>
