magic
tech sky130B
magscale 1 2
timestamp 1683767628
use sky130_fd_pr__hvdfl1sd__example_55959141808278  sky130_fd_pr__hvdfl1sd__example_55959141808278_0
timestamp 1683767628
transform -1 0 0 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 7187394
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7186602
<< end >>
